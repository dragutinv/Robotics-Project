// __  ___ __ ___  _ __   ___  ___ 
// \ \/ / '__/ _ \| '_ \ / _ \/ __|
//  >  <| | | (_) | | | | (_) \__ \
// /_/\_\_|  \___/|_| |_|\___/|___/
// 
// Xronos synthesizer version
// Run date: Tue 17 Nov 2015 18:39:01 +0000
// 

module Generation(Bout_ACK, Rout_COUNT, Rout_SEND, Gin_SEND, Gin_ACK, Bin_ACK, Rout_ACK, Gout_DATA, Rout_DATA, Bout_COUNT, CLK, Gout_RDY, Gout_COUNT, Bin_SEND, Bout_SEND, Gin_DATA, Rin_SEND, Rin_COUNT, Bout_DATA, Bin_COUNT, Gin_COUNT, RESET, Bout_RDY, Bin_DATA, Gout_SEND, Rin_DATA, Rout_RDY, Rin_ACK, Gout_ACK);
input		Bout_ACK;
output	[15:0]	Rout_COUNT;
output		Rout_SEND;
input		Gin_SEND;
output		Gin_ACK;
output		Bin_ACK;
wire		doneCountIm_done;
input		Rout_ACK;
wire		getValueRGB_done;
wire		drawRectangle_done;
output	[7:0]	Gout_DATA;
output	[7:0]	Rout_DATA;
output	[15:0]	Bout_COUNT;
input		CLK;
input		Gout_RDY;
output	[15:0]	Gout_COUNT;
wire		send_go;
input		Bin_SEND;
output		Bout_SEND;
input	[7:0]	Gin_DATA;
wire		doneCountIm_go;
wire		drawRectangle_go;
input		Rin_SEND;
input	[15:0]	Rin_COUNT;
wire		getValueRGB_go;
output	[7:0]	Bout_DATA;
input	[15:0]	Bin_COUNT;
input	[15:0]	Gin_COUNT;
input		RESET;
input		Bout_RDY;
wire		send_done;
input	[7:0]	Bin_DATA;
output		Gout_SEND;
input	[7:0]	Rin_DATA;
input		Rout_RDY;
output		Rin_ACK;
input		Gout_ACK;
wire	[31:0]	bus_0094ee07_;
wire		bus_0063b29b_;
wire		bus_00d78df8_;
wire		bus_00367a8d_;
wire	[7:0]	bus_0044a59b_;
wire	[7:0]	bus_01764bef_;
wire		bus_003c431c_;
wire		bus_00cbefce_;
wire		bus_003a8164_;
wire	[2:0]	bus_01c9832e_;
wire	[31:0]	bus_017e46bf_;
wire	[31:0]	drawRectangle_u269;
wire	[7:0]	drawRectangle_u262;
wire	[2:0]	drawRectangle_u259;
wire	[7:0]	drawRectangle_u258;
wire	[7:0]	drawRectangle_u266;
wire		drawRectangle_u272;
wire	[31:0]	drawRectangle_u261;
wire	[7:0]	drawRectangle_u254;
wire		Generation_drawRectangle_instance_DONE;
wire	[7:0]	drawRectangle_u270;
wire		drawRectangle;
wire	[31:0]	drawRectangle_u273;
wire	[2:0]	drawRectangle_u275;
wire	[31:0]	drawRectangle_u257;
wire	[31:0]	drawRectangle_u253;
wire		drawRectangle_u256;
wire	[2:0]	drawRectangle_u255;
wire	[2:0]	drawRectangle_u267;
wire	[2:0]	drawRectangle_u271;
wire	[2:0]	drawRectangle_u263;
wire		drawRectangle_u268;
wire		drawRectangle_u264;
wire	[31:0]	drawRectangle_u265;
wire	[7:0]	drawRectangle_u274;
wire		drawRectangle_u260;
wire		bus_01530c78_;
wire		getValueRGB_u215;
wire	[2:0]	getValueRGB_u212;
wire	[31:0]	getValueRGB_u198;
wire		getValueRGB_u199;
wire		getValueRGB_u213;
wire		getValueRGB_u201;
wire	[31:0]	getValueRGB_u206;
wire	[2:0]	getValueRGB_u208;
wire	[7:0]	getValueRGB_u207;
wire		getValueRGB;
wire	[31:0]	getValueRGB_u202;
wire		Generation_getValueRGB_instance_DONE;
wire		getValueRGB_u205;
wire	[7:0]	getValueRGB_u211;
wire	[31:0]	getValueRGB_u200;
wire	[7:0]	getValueRGB_u203;
wire	[31:0]	getValueRGB_u210;
wire		getValueRGB_u209;
wire	[2:0]	getValueRGB_u204;
wire		getValueRGB_u214;
wire		bus_00c4eeea_;
wire		bus_01ad823d_;
wire		bus_012df243_;
wire	[7:0]	bus_01dc999c_;
wire		bus_01db46e6_;
wire	[31:0]	doneCountIm_u11;
wire		Generation_doneCountIm_instance_DONE;
wire		doneCountIm;
wire	[2:0]	bus_01fe6336_;
wire		bus_0086d7cf_;
wire	[7:0]	bus_00287f7c_;
wire		bus_0185bd7a_;
wire	[31:0]	bus_01867765_;
wire		bus_0136da55_;
wire		bus_003f9e84_;
wire		bus_01188a3b_;
wire	[7:0]	bus_0072ed28_;
wire		bus_01d34608_;
wire		bus_00f8e3ae_;
wire		bus_01bb2165_;
wire		bus_0042f76c_;
wire	[7:0]	bus_00c1d8fc_;
wire	[2:0]	bus_015b9c7d_;
wire	[7:0]	bus_015536f1_;
wire		bus_007b17d0_;
wire		bus_01d90de5_;
wire	[31:0]	bus_004d0152_;
wire		bus_00dbd379_;
wire		bus_01d5d31c_;
wire	[31:0]	bus_00e65a1a_;
wire		bus_01169eaf_;
wire	[7:0]	bus_005e8953_;
wire		bus_0106a06d_;
wire		bus_01bd7297_;
wire		bus_016bc16f_;
wire	[2:0]	bus_005bc28e_;
wire	[31:0]	bus_01465e99_;
wire		bus_00a84917_;
wire	[7:0]	bus_016572b8_;
wire		bus_0143eb1d_;
wire		bus_01818ac0_;
wire		bus_004cb6d6_;
wire		bus_017f06fa_;
wire		bus_019964a1_;
wire	[7:0]	bus_010ccceb_;
wire	[7:0]	bus_00ac07b4_;
wire	[31:0]	bus_00098098_;
wire		bus_001efe58_;
wire	[2:0]	bus_00e47af6_;
wire		bus_003255c0_;
wire		bus_0159ecfe_;
wire	[2:0]	bus_016e703b_;
wire		bus_015957dd_;
wire	[7:0]	bus_013a971b_;
wire	[31:0]	bus_011fbfd3_;
wire		bus_01d84fc4_;
wire		scheduler_u397;
wire		scheduler_u395;
wire		scheduler;
wire		Generation_scheduler_instance_DONE;
wire		scheduler_u399;
wire		scheduler_u398;
wire		scheduler_u400;
wire		scheduler_u401;
wire		scheduler_u396;
wire		scheduler_u403;
wire		scheduler_u402;
wire		send_u296;
wire	[2:0]	send_u295;
wire	[2:0]	send_u298;
wire	[15:0]	send_u303;
wire	[7:0]	send_u299;
wire		send_u288;
wire	[2:0]	send_u292;
wire		send;
wire	[31:0]	send_u294;
wire	[31:0]	send_u289;
wire		send_u306;
wire		send_u290;
wire		send_u293;
wire	[31:0]	send_u297;
wire	[7:0]	send_u300;
wire	[31:0]	send_u291;
wire		send_u307;
wire	[7:0]	send_u305;
wire	[31:0]	send_u287;
wire	[15:0]	send_u301;
wire	[15:0]	send_u304;
wire		send_u302;
wire		Generation_send_instance_DONE;
assign Rout_COUNT=send_u303;
assign Rout_SEND=send_u306;
assign Gin_ACK=getValueRGB_u215;
assign Bin_ACK=getValueRGB_u213;
assign doneCountIm_done=bus_00a84917_;
assign getValueRGB_done=bus_01169eaf_;
assign drawRectangle_done=bus_01d5d31c_;
assign Gout_DATA=send_u300;
assign Rout_DATA=send_u299;
assign Bout_COUNT=send_u301;
assign Gout_COUNT=send_u304;
assign send_go=scheduler_u401;
assign Bout_SEND=send_u302;
assign doneCountIm_go=scheduler_u402;
assign drawRectangle_go=scheduler_u403;
assign getValueRGB_go=scheduler_u400;
assign Bout_DATA=send_u305;
assign send_done=bus_00f8e3ae_;
assign Gout_SEND=send_u307;
assign Rin_ACK=getValueRGB_u214;
Generation_stateVar_count_x Generation_stateVar_count_x_1(.bus_00236c7e_(CLK), 
  .bus_01a7c757_(bus_01d34608_), .bus_01a0ff1b_(getValueRGB), .bus_01ee5dfb_(getValueRGB_u198), 
  .bus_00d15ba1_(doneCountIm), .bus_01f5fd62_(32'h0), .bus_00a1dfc0_(send), .bus_01dffd60_(send_u287), 
  .bus_0094ee07_(bus_0094ee07_));
Generation_stateVar_state_s1 Generation_stateVar_state_s1_1(.bus_00df16be_(CLK), 
  .bus_004e21ba_(bus_01d34608_), .bus_0081cf58_(scheduler_u396), .bus_013a527d_(scheduler_u397), 
  .bus_0063b29b_(bus_0063b29b_));
Generation_simplememoryreferee_0085b1af_ Generation_simplememoryreferee_0085b1af__1(.bus_009e783e_(CLK), 
  .bus_01e836f8_(bus_01d34608_), .bus_01b0e5fe_(bus_01818ac0_), .bus_012fcde4_(bus_016572b8_), 
  .bus_00133f6a_(getValueRGB_u201), .bus_01276f1b_(getValueRGB_u203), .bus_0010c2f2_(getValueRGB_u202), 
  .bus_00408e3d_(3'h1), .bus_00ca0c9a_(drawRectangle), .bus_00014f14_(8'h0), .bus_012e1581_(drawRectangle_u253), 
  .bus_00822723_(3'h1), .bus_005af008_(send_u290), .bus_01541838_(send_u291), .bus_01371af9_(3'h1), 
  .bus_01764bef_(bus_01764bef_), .bus_017e46bf_(bus_017e46bf_), .bus_003c431c_(bus_003c431c_), 
  .bus_00367a8d_(bus_00367a8d_), .bus_01c9832e_(bus_01c9832e_), .bus_003a8164_(bus_003a8164_), 
  .bus_00d78df8_(bus_00d78df8_), .bus_0044a59b_(bus_0044a59b_), .bus_00cbefce_(bus_00cbefce_));
Generation_drawRectangle Generation_drawRectangle_instance(.CLK(CLK), .RESET(bus_01d34608_), 
  .GO(drawRectangle_go), .port_006e546a_(bus_00d78df8_), .port_01a1bc5b_(bus_0185bd7a_), 
  .port_01ea4bba_(bus_016bc16f_), .port_009296ab_(bus_004cb6d6_), .port_00a4b213_(bus_00dbd379_), 
  .port_004a5ee2_(bus_01d84fc4_), .RESULT(drawRectangle), .RESULT_u1914(drawRectangle_u253), 
  .RESULT_u1915(drawRectangle_u254), .RESULT_u1916(drawRectangle_u255), .RESULT_u1933(drawRectangle_u256), 
  .RESULT_u1934(drawRectangle_u257), .RESULT_u1935(drawRectangle_u258), .RESULT_u1936(drawRectangle_u259), 
  .RESULT_u1921(drawRectangle_u260), .RESULT_u1922(drawRectangle_u261), .RESULT_u1923(drawRectangle_u262), 
  .RESULT_u1924(drawRectangle_u263), .RESULT_u1925(drawRectangle_u264), .RESULT_u1926(drawRectangle_u265), 
  .RESULT_u1927(drawRectangle_u266), .RESULT_u1928(drawRectangle_u267), .RESULT_u1917(drawRectangle_u268), 
  .RESULT_u1918(drawRectangle_u269), .RESULT_u1919(drawRectangle_u270), .RESULT_u1920(drawRectangle_u271), 
  .RESULT_u1929(drawRectangle_u272), .RESULT_u1930(drawRectangle_u273), .RESULT_u1931(drawRectangle_u274), 
  .RESULT_u1932(drawRectangle_u275), .DONE(Generation_drawRectangle_instance_DONE));
Generation_stateVar_state_s0 Generation_stateVar_state_s0_1(.bus_0122c06d_(CLK), 
  .bus_00873bde_(bus_01d34608_), .bus_011920d6_(scheduler), .bus_0020f994_(scheduler_u395), 
  .bus_01530c78_(bus_01530c78_));
Generation_getValueRGB Generation_getValueRGB_instance(.CLK(CLK), .RESET(bus_01d34608_), 
  .GO(getValueRGB_go), .port_007bdc5b_(bus_0094ee07_), .port_01263d81_(bus_00e65a1a_), 
  .port_000d5d4f_(bus_003a8164_), .port_009075e0_(bus_017f06fa_), .port_01f1afae_(bus_01bb2165_), 
  .port_004cc74e_(Gin_DATA), .port_0040ae5e_(Bin_DATA), .port_00960a11_(Rin_DATA), 
  .RESULT(getValueRGB), .RESULT_u1937(getValueRGB_u198), .RESULT_u1938(getValueRGB_u199), 
  .RESULT_u1939(getValueRGB_u200), .RESULT_u1944(getValueRGB_u201), .RESULT_u1945(getValueRGB_u202), 
  .RESULT_u1946(getValueRGB_u203), .RESULT_u1947(getValueRGB_u204), .RESULT_u1948(getValueRGB_u205), 
  .RESULT_u1949(getValueRGB_u206), .RESULT_u1950(getValueRGB_u207), .RESULT_u1951(getValueRGB_u208), 
  .RESULT_u1940(getValueRGB_u209), .RESULT_u1941(getValueRGB_u210), .RESULT_u1942(getValueRGB_u211), 
  .RESULT_u1943(getValueRGB_u212), .RESULT_u1952(getValueRGB_u213), .RESULT_u1953(getValueRGB_u214), 
  .RESULT_u1954(getValueRGB_u215), .DONE(Generation_getValueRGB_instance_DONE));
Generation_Kicker_57 Generation_Kicker_57_1(.CLK(CLK), .RESET(bus_01d34608_), .bus_00c4eeea_(bus_00c4eeea_));
Generation_stateVar_state_s2 Generation_stateVar_state_s2_1(.bus_0168a69b_(CLK), 
  .bus_01920bdc_(bus_01d34608_), .bus_0105be8f_(scheduler_u398), .bus_01b9532b_(scheduler_u399), 
  .bus_01ad823d_(bus_01ad823d_));
Generation_structuralmemory_0156af01_ Generation_structuralmemory_0156af01__1(.CLK_u49(CLK), 
  .bus_0073ced7_(bus_01d34608_), .bus_00fc033f_(bus_00098098_), .bus_00b8b050_(3'h1), 
  .bus_0140811d_(bus_019964a1_), .bus_008c32f9_(bus_003255c0_), .bus_002bf4e6_(bus_00ac07b4_), 
  .bus_00a404ce_(bus_011fbfd3_), .bus_0192694e_(3'h1), .bus_0141e826_(bus_015957dd_), 
  .bus_00d571fa_(8'hff), .bus_01dc999c_(bus_01dc999c_), .bus_01db46e6_(bus_01db46e6_), 
  .bus_012df243_(bus_012df243_));
Generation_doneCountIm Generation_doneCountIm_instance(.CLK(CLK), .RESET(bus_01d34608_), 
  .GO(doneCountIm_go), .RESULT(doneCountIm), .RESULT_u1955(doneCountIm_u11), .DONE(Generation_doneCountIm_instance_DONE));
Generation_simplememoryreferee_000742eb_ Generation_simplememoryreferee_000742eb__1(.bus_0019d89f_(CLK), 
  .bus_00dcc243_(bus_01d34608_), .bus_0057a34a_(bus_0143eb1d_), .bus_013da532_(8'h0), 
  .bus_00660791_(drawRectangle_u256), .bus_007fe65e_(8'h0), .bus_01d1ac5f_(drawRectangle_u257), 
  .bus_01679577_(3'h1), .bus_00287f7c_(bus_00287f7c_), .bus_01867765_(bus_01867765_), 
  .bus_0136da55_(bus_0136da55_), .bus_0086d7cf_(bus_0086d7cf_), .bus_01fe6336_(bus_01fe6336_), 
  .bus_0185bd7a_(bus_0185bd7a_));
Generation_structuralmemory_00c0d3f6_ Generation_structuralmemory_00c0d3f6__1(.CLK_u50(CLK), 
  .bus_01d2754e_(bus_01d34608_), .bus_000dbf39_(bus_004d0152_), .bus_0149775b_(3'h1), 
  .bus_003a8ec4_(bus_0042f76c_), .bus_01674500_(bus_01d90de5_), .bus_0108036b_(bus_015536f1_), 
  .bus_01ae55ef_(bus_01465e99_), .bus_00a5d728_(3'h1), .bus_01563c6d_(bus_01bd7297_), 
  .bus_000f6b16_(8'h0), .bus_0072ed28_(bus_0072ed28_), .bus_01188a3b_(bus_01188a3b_), 
  .bus_003f9e84_(bus_003f9e84_));
Generation_globalreset_physical_018187f8_ Generation_globalreset_physical_018187f8__1(.bus_00cbf5a7_(CLK), 
  .bus_0058fdd8_(RESET), .bus_01d34608_(bus_01d34608_));
assign bus_00f8e3ae_=Generation_send_instance_DONE&{1{Generation_send_instance_DONE}};
Generation_simplememoryreferee_0062bad9_ Generation_simplememoryreferee_0062bad9__1(.bus_006120d5_(CLK), 
  .bus_00b2b57c_(bus_01d34608_), .bus_018943bd_(bus_01188a3b_), .bus_007f922a_(bus_0072ed28_), 
  .bus_0128b244_(getValueRGB_u209), .bus_01da6bec_(getValueRGB_u211), .bus_00a675df_(getValueRGB_u210), 
  .bus_00b36d07_(3'h1), .bus_011ac12c_(drawRectangle_u268), .bus_004c87c7_(8'h0), 
  .bus_01fc3728_(drawRectangle_u269), .bus_005db036_(3'h1), .bus_01966503_(send_u293), 
  .bus_005f1004_(send_u294), .bus_00837cdf_(3'h1), .bus_015536f1_(bus_015536f1_), 
  .bus_004d0152_(bus_004d0152_), .bus_01d90de5_(bus_01d90de5_), .bus_0042f76c_(bus_0042f76c_), 
  .bus_015b9c7d_(bus_015b9c7d_), .bus_01bb2165_(bus_01bb2165_), .bus_00dbd379_(bus_00dbd379_), 
  .bus_00c1d8fc_(bus_00c1d8fc_), .bus_007b17d0_(bus_007b17d0_));
assign bus_01d5d31c_=Generation_drawRectangle_instance_DONE&{1{Generation_drawRectangle_instance_DONE}};
Generation_stateVar_count_y Generation_stateVar_count_y_1(.bus_0168294f_(CLK), 
  .bus_017039a6_(bus_01d34608_), .bus_0130359b_(getValueRGB_u199), .bus_00d547ca_(getValueRGB_u200), 
  .bus_007d4ec1_(send_u288), .bus_00272892_(send_u289), .bus_00e65a1a_(bus_00e65a1a_));
assign bus_01169eaf_=Generation_getValueRGB_instance_DONE&{1{Generation_getValueRGB_instance_DONE}};
Generation_simplememoryreferee_01801ae8_ Generation_simplememoryreferee_01801ae8__1(.bus_005cefdf_(CLK), 
  .bus_01883661_(bus_01d34608_), .bus_01533ec6_(bus_003f9e84_), .bus_01625b66_(8'h0), 
  .bus_005222c2_(drawRectangle_u260), .bus_004e4c93_(8'h0), .bus_008195d8_(drawRectangle_u261), 
  .bus_0133852a_(3'h1), .bus_005e8953_(bus_005e8953_), .bus_01465e99_(bus_01465e99_), 
  .bus_01bd7297_(bus_01bd7297_), .bus_0106a06d_(bus_0106a06d_), .bus_005bc28e_(bus_005bc28e_), 
  .bus_016bc16f_(bus_016bc16f_));
assign bus_00a84917_=Generation_doneCountIm_instance_DONE&{1{Generation_doneCountIm_instance_DONE}};
Generation_structuralmemory_01173ea4_ Generation_structuralmemory_01173ea4__1(.CLK_u51(CLK), 
  .bus_00145df3_(bus_01d34608_), .bus_012e52ce_(bus_017e46bf_), .bus_0040491c_(3'h1), 
  .bus_005d0e89_(bus_00367a8d_), .bus_0041c93d_(bus_003c431c_), .bus_00133706_(bus_01764bef_), 
  .bus_0085d248_(bus_01867765_), .bus_00aaeacd_(3'h1), .bus_01b5bcf2_(bus_0136da55_), 
  .bus_00bb37ab_(8'h0), .bus_016572b8_(bus_016572b8_), .bus_01818ac0_(bus_01818ac0_), 
  .bus_0143eb1d_(bus_0143eb1d_));
Generation_simplememoryreferee_0173d745_ Generation_simplememoryreferee_0173d745__1(.bus_00527630_(CLK), 
  .bus_01cd82ec_(bus_01d34608_), .bus_01248bfe_(bus_01db46e6_), .bus_005611d2_(bus_01dc999c_), 
  .bus_00769b40_(getValueRGB_u205), .bus_0149134b_(getValueRGB_u207), .bus_0149fcb3_(getValueRGB_u206), 
  .bus_0148efea_(3'h1), .bus_0018bf4d_(drawRectangle_u264), .bus_006f81ca_(8'hff), 
  .bus_014b9e03_(drawRectangle_u265), .bus_0065e7ab_(3'h1), .bus_00309326_(send_u296), 
  .bus_01835b38_(send_u297), .bus_01b43d37_(3'h1), .bus_00ac07b4_(bus_00ac07b4_), 
  .bus_00098098_(bus_00098098_), .bus_003255c0_(bus_003255c0_), .bus_019964a1_(bus_019964a1_), 
  .bus_00e47af6_(bus_00e47af6_), .bus_017f06fa_(bus_017f06fa_), .bus_004cb6d6_(bus_004cb6d6_), 
  .bus_010ccceb_(bus_010ccceb_), .bus_001efe58_(bus_001efe58_));
Generation_simplememoryreferee_00377ebe_ Generation_simplememoryreferee_00377ebe__1(.bus_014779db_(CLK), 
  .bus_01911ea6_(bus_01d34608_), .bus_019e8d0b_(bus_012df243_), .bus_00efbc69_(8'h0), 
  .bus_004c6569_(drawRectangle_u272), .bus_007ef2a5_(8'hff), .bus_00d7d56a_(drawRectangle_u273), 
  .bus_0033b983_(3'h1), .bus_013a971b_(bus_013a971b_), .bus_011fbfd3_(bus_011fbfd3_), 
  .bus_015957dd_(bus_015957dd_), .bus_0159ecfe_(bus_0159ecfe_), .bus_016e703b_(bus_016e703b_), 
  .bus_01d84fc4_(bus_01d84fc4_));
Generation_scheduler Generation_scheduler_instance(.CLK(CLK), .RESET(bus_01d34608_), 
  .GO(bus_00c4eeea_), .port_0032333f_(bus_01530c78_), .port_01ce98f6_(bus_0063b29b_), 
  .port_00c47705_(bus_01ad823d_), .port_00dad65c_(bus_0094ee07_), .port_012c5997_(doneCountIm_done), 
  .port_00a666cf_(Rin_SEND), .port_001c856e_(Rout_RDY), .port_000be277_(Gout_RDY), 
  .port_012fe075_(getValueRGB_done), .port_00429cca_(send_done), .port_00d4319a_(Bout_RDY), 
  .port_00c133f5_(Gin_SEND), .port_010c32d0_(drawRectangle_done), .port_01d1c7ea_(Bin_SEND), 
  .RESULT(scheduler), .RESULT_u1956(scheduler_u395), .RESULT_u1957(scheduler_u396), 
  .RESULT_u1958(scheduler_u397), .RESULT_u1959(scheduler_u398), .RESULT_u1960(scheduler_u399), 
  .RESULT_u1961(scheduler_u400), .RESULT_u1962(scheduler_u401), .RESULT_u1964(scheduler_u402), 
  .RESULT_u1963(scheduler_u403), .DONE(Generation_scheduler_instance_DONE));
Generation_send Generation_send_instance(.CLK(CLK), .RESET(bus_01d34608_), .GO(send_go), 
  .port_00bf371b_(bus_0094ee07_), .port_0158b5cb_(bus_00e65a1a_), .port_00f76336_(bus_00cbefce_), 
  .port_006cd08b_(bus_0044a59b_), .port_00b84c6a_(bus_007b17d0_), .port_01177a51_(bus_00c1d8fc_), 
  .port_0197dc98_(bus_001efe58_), .port_0079b3b6_(bus_010ccceb_), .RESULT(send), 
  .RESULT_u1965(send_u287), .RESULT_u1966(send_u288), .RESULT_u1967(send_u289), 
  .RESULT_u1971(send_u290), .RESULT_u1972(send_u291), .RESULT_u1973(send_u292), 
  .RESULT_u1968(send_u293), .RESULT_u1969(send_u294), .RESULT_u1970(send_u295), 
  .RESULT_u1974(send_u296), .RESULT_u1975(send_u297), .RESULT_u1976(send_u298), 
  .RESULT_u1979(send_u299), .RESULT_u1978(send_u300), .RESULT_u1977(send_u301), 
  .RESULT_u1980(send_u302), .RESULT_u1981(send_u303), .RESULT_u1983(send_u304), 
  .RESULT_u1982(send_u305), .RESULT_u1984(send_u306), .RESULT_u1985(send_u307), 
  .DONE(Generation_send_instance_DONE));
endmodule



module Generation_endianswapper_00cebe92_(endianswapper_00cebe92_in, endianswapper_00cebe92_out);
input	[31:0]	endianswapper_00cebe92_in;
output	[31:0]	endianswapper_00cebe92_out;
assign endianswapper_00cebe92_out=endianswapper_00cebe92_in;
endmodule



module Generation_endianswapper_0107c13c_(endianswapper_0107c13c_in, endianswapper_0107c13c_out);
input	[31:0]	endianswapper_0107c13c_in;
output	[31:0]	endianswapper_0107c13c_out;
assign endianswapper_0107c13c_out=endianswapper_0107c13c_in;
endmodule



module Generation_stateVar_count_x(bus_00236c7e_, bus_01a7c757_, bus_01a0ff1b_, bus_01ee5dfb_, bus_00d15ba1_, bus_01f5fd62_, bus_00a1dfc0_, bus_01dffd60_, bus_0094ee07_);
input		bus_00236c7e_;
input		bus_01a7c757_;
input		bus_01a0ff1b_;
input	[31:0]	bus_01ee5dfb_;
input		bus_00d15ba1_;
input	[31:0]	bus_01f5fd62_;
input		bus_00a1dfc0_;
input	[31:0]	bus_01dffd60_;
output	[31:0]	bus_0094ee07_;
wire		or_00d7d677_u0;
wire	[31:0]	mux_018c344f_u0;
wire	[31:0]	endianswapper_00cebe92_out;
wire	[31:0]	endianswapper_0107c13c_out;
reg	[31:0]	stateVar_count_x_u11=32'h0;
assign or_00d7d677_u0=bus_01a0ff1b_|bus_00d15ba1_|bus_00a1dfc0_;
assign mux_018c344f_u0=({32{bus_01a0ff1b_}}&bus_01ee5dfb_)|({32{bus_00d15ba1_}}&32'h0)|({32{bus_00a1dfc0_}}&bus_01dffd60_);
Generation_endianswapper_00cebe92_ Generation_endianswapper_00cebe92__1(.endianswapper_00cebe92_in(mux_018c344f_u0), 
  .endianswapper_00cebe92_out(endianswapper_00cebe92_out));
Generation_endianswapper_0107c13c_ Generation_endianswapper_0107c13c__1(.endianswapper_0107c13c_in(stateVar_count_x_u11), 
  .endianswapper_0107c13c_out(endianswapper_0107c13c_out));
always @(posedge bus_00236c7e_ or posedge bus_01a7c757_)
begin
if (bus_01a7c757_)
stateVar_count_x_u11<=32'h0;
else if (or_00d7d677_u0)
stateVar_count_x_u11<=endianswapper_00cebe92_out;
end
assign bus_0094ee07_=endianswapper_0107c13c_out;
endmodule



module Generation_stateVar_state_s1(bus_00df16be_, bus_004e21ba_, bus_0081cf58_, bus_013a527d_, bus_0063b29b_);
input		bus_00df16be_;
input		bus_004e21ba_;
input		bus_0081cf58_;
input		bus_013a527d_;
output		bus_0063b29b_;
reg		stateVar_state_s1_u34=1'h0;
assign bus_0063b29b_=stateVar_state_s1_u34;
always @(posedge bus_00df16be_ or posedge bus_004e21ba_)
begin
if (bus_004e21ba_)
stateVar_state_s1_u34<=1'h0;
else if (bus_0081cf58_)
stateVar_state_s1_u34<=bus_013a527d_;
end
endmodule



module Generation_simplememoryreferee_0085b1af_(bus_009e783e_, bus_01e836f8_, bus_01b0e5fe_, bus_012fcde4_, bus_00133f6a_, bus_01276f1b_, bus_0010c2f2_, bus_00408e3d_, bus_00ca0c9a_, bus_00014f14_, bus_012e1581_, bus_00822723_, bus_005af008_, bus_01541838_, bus_01371af9_, bus_01764bef_, bus_017e46bf_, bus_003c431c_, bus_00367a8d_, bus_01c9832e_, bus_003a8164_, bus_00d78df8_, bus_0044a59b_, bus_00cbefce_);
input		bus_009e783e_;
input		bus_01e836f8_;
input		bus_01b0e5fe_;
input	[7:0]	bus_012fcde4_;
input		bus_00133f6a_;
input	[7:0]	bus_01276f1b_;
input	[31:0]	bus_0010c2f2_;
input	[2:0]	bus_00408e3d_;
input		bus_00ca0c9a_;
input	[7:0]	bus_00014f14_;
input	[31:0]	bus_012e1581_;
input	[2:0]	bus_00822723_;
input		bus_005af008_;
input	[31:0]	bus_01541838_;
input	[2:0]	bus_01371af9_;
output	[7:0]	bus_01764bef_;
output	[31:0]	bus_017e46bf_;
output		bus_003c431c_;
output		bus_00367a8d_;
output	[2:0]	bus_01c9832e_;
output		bus_003a8164_;
output		bus_00d78df8_;
output	[7:0]	bus_0044a59b_;
output		bus_00cbefce_;
wire		and_01b62546_u0;
reg		done_qual_u147=1'h0;
wire		or_0042eabf_u0;
wire		not_00209fed_u0;
wire		or_01805839_u0;
wire		or_01d0e7e1_u0;
wire	[7:0]	mux_0092760b_u0;
wire		not_00729a48_u0;
wire		and_00148a93_u0;
wire		or_009d019e_u0;
wire		and_00953dcf_u0;
reg		done_qual_u148_u0=1'h0;
wire	[31:0]	mux_00f089f3_u0;
reg		done_qual_u149_u0=1'h0;
wire		not_0089f43a_u0;
wire		or_018e20f5_u0;
assign and_01b62546_u0=or_009d019e_u0&bus_01b0e5fe_;
always @(posedge bus_009e783e_)
begin
if (bus_01e836f8_)
done_qual_u147<=1'h0;
else done_qual_u147<=bus_00ca0c9a_;
end
assign or_0042eabf_u0=bus_00133f6a_|done_qual_u148_u0;
assign not_00209fed_u0=~bus_01b0e5fe_;
assign or_01805839_u0=bus_005af008_|done_qual_u149_u0;
assign or_01d0e7e1_u0=bus_00133f6a_|bus_00ca0c9a_;
assign bus_01764bef_=mux_0092760b_u0;
assign bus_017e46bf_=mux_00f089f3_u0;
assign bus_003c431c_=or_01d0e7e1_u0;
assign bus_00367a8d_=or_018e20f5_u0;
assign bus_01c9832e_=3'h1;
assign bus_003a8164_=and_00148a93_u0;
assign bus_00d78df8_=and_01b62546_u0;
assign bus_0044a59b_=bus_012fcde4_;
assign bus_00cbefce_=and_00953dcf_u0;
assign mux_0092760b_u0=(bus_00133f6a_)?bus_01276f1b_:8'h0;
assign not_00729a48_u0=~bus_01b0e5fe_;
assign and_00148a93_u0=or_0042eabf_u0&bus_01b0e5fe_;
assign or_009d019e_u0=bus_00ca0c9a_|done_qual_u147;
assign and_00953dcf_u0=or_01805839_u0&bus_01b0e5fe_;
always @(posedge bus_009e783e_)
begin
if (bus_01e836f8_)
done_qual_u148_u0<=1'h0;
else done_qual_u148_u0<=bus_00133f6a_;
end
assign mux_00f089f3_u0=({32{bus_00133f6a_}}&bus_0010c2f2_)|({32{bus_00ca0c9a_}}&bus_012e1581_)|({32{bus_005af008_}}&bus_01541838_);
always @(posedge bus_009e783e_)
begin
if (bus_01e836f8_)
done_qual_u149_u0<=1'h0;
else done_qual_u149_u0<=bus_005af008_;
end
assign not_0089f43a_u0=~bus_01b0e5fe_;
assign or_018e20f5_u0=bus_00133f6a_|bus_00ca0c9a_|bus_005af008_;
endmodule



module Generation_drawRectangle(CLK, RESET, GO, port_006e546a_, port_00a4b213_, port_01ea4bba_, port_009296ab_, port_004a5ee2_, port_01a1bc5b_, RESULT, RESULT_u1914, RESULT_u1915, RESULT_u1916, RESULT_u1917, RESULT_u1918, RESULT_u1919, RESULT_u1920, RESULT_u1921, RESULT_u1922, RESULT_u1923, RESULT_u1924, RESULT_u1925, RESULT_u1926, RESULT_u1927, RESULT_u1928, RESULT_u1929, RESULT_u1930, RESULT_u1931, RESULT_u1932, RESULT_u1933, RESULT_u1934, RESULT_u1935, RESULT_u1936, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_006e546a_;
input		port_00a4b213_;
input		port_01ea4bba_;
input		port_009296ab_;
input		port_004a5ee2_;
input		port_01a1bc5b_;
output		RESULT;
output	[31:0]	RESULT_u1914;
output	[7:0]	RESULT_u1915;
output	[2:0]	RESULT_u1916;
output		RESULT_u1917;
output	[31:0]	RESULT_u1918;
output	[7:0]	RESULT_u1919;
output	[2:0]	RESULT_u1920;
output		RESULT_u1921;
output	[31:0]	RESULT_u1922;
output	[7:0]	RESULT_u1923;
output	[2:0]	RESULT_u1924;
output		RESULT_u1925;
output	[31:0]	RESULT_u1926;
output	[7:0]	RESULT_u1927;
output	[2:0]	RESULT_u1928;
output		RESULT_u1929;
output	[31:0]	RESULT_u1930;
output	[7:0]	RESULT_u1931;
output	[2:0]	RESULT_u1932;
output		RESULT_u1933;
output	[31:0]	RESULT_u1934;
output	[7:0]	RESULT_u1935;
output	[2:0]	RESULT_u1936;
output		DONE;
wire	[31:0]	add;
wire	[31:0]	add_u1105;
wire		and_u2609_u0;
wire		or_u715_u0;
reg		reg_0169ebdc_u0=1'h0;
wire	[31:0]	add_u1106;
wire	[31:0]	add_u1107;
wire		or_u716_u0;
reg		reg_00f6950d_u0=1'h0;
wire		and_u2610_u0;
wire	[31:0]	add_u1108;
wire	[31:0]	add_u1109;
wire		or_u717_u0;
wire		and_u2611_u0;
reg		reg_01e67662_u0=1'h0;
wire	[31:0]	add_u1110;
wire	[31:0]	add_u1111;
wire		and_u2612_u0;
reg		reg_01c4e2a8_u0=1'h0;
wire		or_u718_u0;
wire	[31:0]	add_u1112;
wire	[31:0]	add_u1113;
wire		and_u2613_u0;
reg		reg_01e2c2e3_u0=1'h0;
wire		or_u719_u0;
wire	[31:0]	add_u1114;
wire	[31:0]	add_u1115;
wire		and_u2614_u0;
wire		or_u720_u0;
reg		reg_01853ac8_u0=1'h0;
wire	[31:0]	add_u1116;
reg		block_GO_delayed_u40=1'h0;
reg	[31:0]	syncEnable_u351=32'h0;
reg	[31:0]	syncEnable_u352_u0=32'h0;
reg	[31:0]	syncEnable_u353_u0=32'h0;
reg	[31:0]	syncEnable_u354_u0=32'h0;
reg	[31:0]	syncEnable_u355_u0=32'h0;
reg	[31:0]	syncEnable_u356_u0=32'h0;
reg		block_GO_delayed_result_delayed_u6=1'h0;
reg	[31:0]	syncEnable_u357_u0=32'h0;
wire		and_u2615_u0;
wire signed	[31:0]	lessThanEqualTo_b_signed;
wire signed	[31:0]	lessThanEqualTo_a_signed;
wire		lessThanEqualTo;
wire		and_u2616_u0;
wire		not_u547_u0;
wire		and_u2617_u0;
wire		and_u2618_u0;
reg		reg_0016dba7_u0=1'h0;
reg		and_delayed_u62=1'h0;
reg		and_delayed_result_delayed_u10=1'h0;
wire	[31:0]	mux_u486;
reg	[6:0]	latch_01d3911a_reg=7'h0;
wire	[31:0]	latch_01d3911a_out;
wire		or_u721_u0;
wire		and_u2619_u0;
reg		and_delayed_u63_u0=1'h0;
wire	[31:0]	add_u1117;
wire	[31:0]	add_u1118;
wire	[31:0]	add_u1119;
wire	[31:0]	add_u1120;
wire		and_u2620_u0;
reg		reg_009152c6_u0=1'h0;
wire		or_u722_u0;
wire	[31:0]	add_u1121;
wire	[31:0]	add_u1122;
wire	[31:0]	add_u1123;
wire	[31:0]	add_u1124;
wire		or_u723_u0;
wire		and_u2621_u0;
reg		reg_014e0cca_u0=1'h0;
wire	[31:0]	add_u1125;
wire	[31:0]	add_u1126;
wire	[31:0]	add_u1127;
wire	[31:0]	add_u1128;
wire		and_u2622_u0;
wire		or_u724_u0;
reg		reg_008df4c9_u0=1'h0;
wire	[31:0]	add_u1129;
wire	[31:0]	add_u1130;
wire	[31:0]	add_u1131;
wire	[31:0]	add_u1132;
wire		or_u725_u0;
wire		and_u2623_u0;
reg		reg_015b2ecc_u0=1'h0;
wire	[31:0]	add_u1133;
wire	[31:0]	add_u1134;
wire	[31:0]	add_u1135;
wire	[31:0]	add_u1136;
wire		or_u726_u0;
reg		reg_01144fd1_u0=1'h0;
wire		and_u2624_u0;
wire	[31:0]	add_u1137;
wire	[31:0]	add_u1138;
wire	[31:0]	add_u1139;
wire	[31:0]	add_u1140;
reg		reg_0114ad74_u0=1'h0;
wire		and_u2625_u0;
wire		or_u727_u0;
wire	[31:0]	add_u1141;
reg	[31:0]	syncEnable_u358_u0=32'h0;
reg	[31:0]	syncEnable_u359_u0=32'h0;
reg	[31:0]	syncEnable_u360_u0=32'h0;
reg		block_GO_delayed_u41_u0=1'h0;
reg	[31:0]	syncEnable_u361_u0=32'h0;
reg	[31:0]	syncEnable_u362_u0=32'h0;
reg		block_GO_delayed_result_delayed_u7_u0=1'h0;
reg	[31:0]	syncEnable_u363_u0=32'h0;
reg	[31:0]	syncEnable_u364_u0=32'h0;
reg		reg_01cf1df3_u0=1'h0;
wire signed	[31:0]	lessThanEqualTo_u11_a_signed;
wire		lessThanEqualTo_u11;
wire signed	[31:0]	lessThanEqualTo_u11_b_signed;
wire		not_u548_u0;
wire		and_u2626_u0;
wire		and_u2627_u0;
reg		and_delayed_result_delayed_u11_u0=1'h0;
wire		and_u2628_u0;
wire	[31:0]	latch_01b87821_out;
reg	[5:0]	latch_01b87821_reg=6'h0;
wire	[31:0]	latch_006cd68c_out;
reg	[6:0]	latch_006cd68c_reg=7'h0;
wire	[31:0]	mux_u487_u0;
wire	[31:0]	latch_0083bde1_out;
reg	[6:0]	latch_0083bde1_reg=7'h0;
wire		or_u728_u0;
wire	[31:0]	mux_u488_u0;
wire		or_u729_u0;
wire		or_u730_u0;
wire	[31:0]	mux_u489_u0;
wire		or_u731_u0;
wire	[31:0]	mux_u490_u0;
reg		reg_017046c7_u0=1'h0;
wire	[31:0]	mux_u491_u0;
wire		or_u732_u0;
wire		or_u733_u0;
wire	[31:0]	mux_u492_u0;
wire		or_u734_u0;
wire	[31:0]	mux_u493_u0;
assign add=32'h1130+mux_u486;
assign add_u1105=32'h0+add;
assign and_u2609_u0=reg_0169ebdc_u0&port_009296ab_;
assign or_u715_u0=and_u2609_u0|RESET;
always @(posedge CLK or posedge block_GO_delayed_u40 or posedge or_u715_u0)
begin
if (or_u715_u0)
reg_0169ebdc_u0<=1'h0;
else if (block_GO_delayed_u40)
reg_0169ebdc_u0<=1'h1;
else reg_0169ebdc_u0<=reg_0169ebdc_u0;
end
assign add_u1106=32'h1130+mux_u486;
assign add_u1107=32'h0+add_u1106;
assign or_u716_u0=and_u2610_u0|RESET;
always @(posedge CLK or posedge block_GO_delayed_u40 or posedge or_u716_u0)
begin
if (or_u716_u0)
reg_00f6950d_u0<=1'h0;
else if (block_GO_delayed_u40)
reg_00f6950d_u0<=1'h1;
else reg_00f6950d_u0<=reg_00f6950d_u0;
end
assign and_u2610_u0=reg_00f6950d_u0&port_006e546a_;
assign add_u1108=32'h1130+mux_u486;
assign add_u1109=32'h0+add_u1108;
assign or_u717_u0=and_u2611_u0|RESET;
assign and_u2611_u0=reg_01e67662_u0&port_00a4b213_;
always @(posedge CLK or posedge block_GO_delayed_u40 or posedge or_u717_u0)
begin
if (or_u717_u0)
reg_01e67662_u0<=1'h0;
else if (block_GO_delayed_u40)
reg_01e67662_u0<=1'h1;
else reg_01e67662_u0<=reg_01e67662_u0;
end
assign add_u1110=32'h25d0+mux_u486;
assign add_u1111=32'h0+add_u1110;
assign and_u2612_u0=reg_01c4e2a8_u0&port_004a5ee2_;
always @(posedge CLK or posedge block_GO_delayed_result_delayed_u6 or posedge or_u718_u0)
begin
if (or_u718_u0)
reg_01c4e2a8_u0<=1'h0;
else if (block_GO_delayed_result_delayed_u6)
reg_01c4e2a8_u0<=1'h1;
else reg_01c4e2a8_u0<=reg_01c4e2a8_u0;
end
assign or_u718_u0=and_u2612_u0|RESET;
assign add_u1112=32'h25d0+mux_u486;
assign add_u1113=32'h0+add_u1112;
assign and_u2613_u0=reg_01e2c2e3_u0&port_01a1bc5b_;
always @(posedge CLK or posedge block_GO_delayed_result_delayed_u6 or posedge or_u719_u0)
begin
if (or_u719_u0)
reg_01e2c2e3_u0<=1'h0;
else if (block_GO_delayed_result_delayed_u6)
reg_01e2c2e3_u0<=1'h1;
else reg_01e2c2e3_u0<=reg_01e2c2e3_u0;
end
assign or_u719_u0=and_u2613_u0|RESET;
assign add_u1114=32'h25d0+mux_u486;
assign add_u1115=32'h0+add_u1114;
assign and_u2614_u0=reg_01853ac8_u0&port_01ea4bba_;
assign or_u720_u0=and_u2614_u0|RESET;
always @(posedge CLK or posedge block_GO_delayed_result_delayed_u6 or posedge or_u720_u0)
begin
if (or_u720_u0)
reg_01853ac8_u0<=1'h0;
else if (block_GO_delayed_result_delayed_u6)
reg_01853ac8_u0<=1'h1;
else reg_01853ac8_u0<=reg_01853ac8_u0;
end
assign add_u1116=mux_u486+32'h1;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u40<=1'h0;
else block_GO_delayed_u40<=and_u2615_u0;
end
always @(posedge CLK)
begin
if (and_u2615_u0)
syncEnable_u351<=add_u1116;
end
always @(posedge CLK)
begin
if (and_u2615_u0)
syncEnable_u352_u0<=add_u1115;
end
always @(posedge CLK)
begin
if (and_u2615_u0)
syncEnable_u353_u0<=add_u1109;
end
always @(posedge CLK)
begin
if (and_u2615_u0)
syncEnable_u354_u0<=add_u1111;
end
always @(posedge CLK)
begin
if (and_u2615_u0)
syncEnable_u355_u0<=add_u1107;
end
always @(posedge CLK)
begin
if (and_u2615_u0)
syncEnable_u356_u0<=add_u1113;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_result_delayed_u6<=1'h0;
else block_GO_delayed_result_delayed_u6<=block_GO_delayed_u40;
end
always @(posedge CLK)
begin
if (and_u2615_u0)
syncEnable_u357_u0<=add_u1105;
end
assign and_u2615_u0=and_u2617_u0&or_u721_u0;
assign lessThanEqualTo_a_signed=mux_u486;
assign lessThanEqualTo_b_signed=32'h32;
assign lessThanEqualTo=lessThanEqualTo_a_signed<=lessThanEqualTo_b_signed;
assign and_u2616_u0=or_u721_u0&not_u547_u0;
assign not_u547_u0=~lessThanEqualTo;
assign and_u2617_u0=or_u721_u0&lessThanEqualTo;
assign and_u2618_u0=and_u2616_u0&or_u721_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0016dba7_u0<=1'h0;
else reg_0016dba7_u0<=and_delayed_result_delayed_u10;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u62<=1'h0;
else and_delayed_u62<=and_u2615_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_u10<=1'h0;
else and_delayed_result_delayed_u10<=and_delayed_u62;
end
assign mux_u486=(reg_0016dba7_u0)?syncEnable_u351:32'h1e;
always @(posedge CLK)
begin
if (reg_017046c7_u0)
latch_01d3911a_reg<=7'h32;
end
assign latch_01d3911a_out=(reg_017046c7_u0)?32'h32:32'h32;
assign or_u721_u0=reg_0016dba7_u0|reg_017046c7_u0;
assign and_u2619_u0=and_u2626_u0&or_u728_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u63_u0<=1'h0;
else and_delayed_u63_u0<=and_u2619_u0;
end
assign add_u1117={mux_u487_u0[24:0], 7'b0}+{mux_u487_u0[26:0], 5'b0};
assign add_u1118={add_u1117[31:5], 5'b0}+{mux_u487_u0[27:0], 4'b0};
assign add_u1119={add_u1118[31:4], 4'b0}+32'h1e;
assign add_u1120=32'h0+{add_u1119[31:4], 4'b1110};
assign and_u2620_u0=reg_009152c6_u0&port_009296ab_;
always @(posedge CLK or posedge block_GO_delayed_u41_u0 or posedge or_u722_u0)
begin
if (or_u722_u0)
reg_009152c6_u0<=1'h0;
else if (block_GO_delayed_u41_u0)
reg_009152c6_u0<=1'h1;
else reg_009152c6_u0<=reg_009152c6_u0;
end
assign or_u722_u0=and_u2620_u0|RESET;
assign add_u1121={mux_u487_u0[24:0], 7'b0}+{mux_u487_u0[26:0], 5'b0};
assign add_u1122={add_u1121[31:5], 5'b0}+{mux_u487_u0[27:0], 4'b0};
assign add_u1123={add_u1122[31:4], 4'b0}+32'h1e;
assign add_u1124=32'h0+{add_u1123[31:4], 4'b1110};
assign or_u723_u0=and_u2621_u0|RESET;
assign and_u2621_u0=reg_014e0cca_u0&port_006e546a_;
always @(posedge CLK or posedge block_GO_delayed_u41_u0 or posedge or_u723_u0)
begin
if (or_u723_u0)
reg_014e0cca_u0<=1'h0;
else if (block_GO_delayed_u41_u0)
reg_014e0cca_u0<=1'h1;
else reg_014e0cca_u0<=reg_014e0cca_u0;
end
assign add_u1125={mux_u487_u0[24:0], 7'b0}+{mux_u487_u0[26:0], 5'b0};
assign add_u1126={add_u1125[31:5], 5'b0}+{mux_u487_u0[27:0], 4'b0};
assign add_u1127={add_u1126[31:4], 4'b0}+32'h1e;
assign add_u1128=32'h0+{add_u1127[31:4], 4'b1110};
assign and_u2622_u0=reg_008df4c9_u0&port_00a4b213_;
assign or_u724_u0=and_u2622_u0|RESET;
always @(posedge CLK or posedge block_GO_delayed_u41_u0 or posedge or_u724_u0)
begin
if (or_u724_u0)
reg_008df4c9_u0<=1'h0;
else if (block_GO_delayed_u41_u0)
reg_008df4c9_u0<=1'h1;
else reg_008df4c9_u0<=reg_008df4c9_u0;
end
assign add_u1129={mux_u487_u0[24:0], 7'b0}+{mux_u487_u0[26:0], 5'b0};
assign add_u1130={add_u1129[31:5], 5'b0}+{mux_u487_u0[27:0], 4'b0};
assign add_u1131={add_u1130[31:4], 4'b0}+32'h32;
assign add_u1132=32'h0+{add_u1131[31:4], 4'b10};
assign or_u725_u0=and_u2623_u0|RESET;
assign and_u2623_u0=reg_015b2ecc_u0&port_004a5ee2_;
always @(posedge CLK or posedge block_GO_delayed_result_delayed_u7_u0 or posedge or_u725_u0)
begin
if (or_u725_u0)
reg_015b2ecc_u0<=1'h0;
else if (block_GO_delayed_result_delayed_u7_u0)
reg_015b2ecc_u0<=1'h1;
else reg_015b2ecc_u0<=reg_015b2ecc_u0;
end
assign add_u1133={mux_u487_u0[24:0], 7'b0}+{mux_u487_u0[26:0], 5'b0};
assign add_u1134={add_u1133[31:5], 5'b0}+{mux_u487_u0[27:0], 4'b0};
assign add_u1135={add_u1134[31:4], 4'b0}+32'h32;
assign add_u1136=32'h0+{add_u1135[31:4], 4'b10};
assign or_u726_u0=and_u2624_u0|RESET;
always @(posedge CLK or posedge block_GO_delayed_result_delayed_u7_u0 or posedge or_u726_u0)
begin
if (or_u726_u0)
reg_01144fd1_u0<=1'h0;
else if (block_GO_delayed_result_delayed_u7_u0)
reg_01144fd1_u0<=1'h1;
else reg_01144fd1_u0<=reg_01144fd1_u0;
end
assign and_u2624_u0=reg_01144fd1_u0&port_01a1bc5b_;
assign add_u1137={mux_u487_u0[24:0], 7'b0}+{mux_u487_u0[26:0], 5'b0};
assign add_u1138={add_u1137[31:5], 5'b0}+{mux_u487_u0[27:0], 4'b0};
assign add_u1139={add_u1138[31:4], 4'b0}+32'h32;
assign add_u1140=32'h0+{add_u1139[31:4], 4'b10};
always @(posedge CLK or posedge block_GO_delayed_result_delayed_u7_u0 or posedge or_u727_u0)
begin
if (or_u727_u0)
reg_0114ad74_u0<=1'h0;
else if (block_GO_delayed_result_delayed_u7_u0)
reg_0114ad74_u0<=1'h1;
else reg_0114ad74_u0<=reg_0114ad74_u0;
end
assign and_u2625_u0=reg_0114ad74_u0&port_01ea4bba_;
assign or_u727_u0=and_u2625_u0|RESET;
assign add_u1141=mux_u487_u0+32'h1;
always @(posedge CLK)
begin
if (and_u2619_u0)
syncEnable_u358_u0<={add_u1120[31:4], 4'b1110};
end
always @(posedge CLK)
begin
if (and_u2619_u0)
syncEnable_u359_u0<={add_u1140[31:4], 4'b10};
end
always @(posedge CLK)
begin
if (and_u2619_u0)
syncEnable_u360_u0<=add_u1141;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u41_u0<=1'h0;
else block_GO_delayed_u41_u0<=and_u2619_u0;
end
always @(posedge CLK)
begin
if (and_u2619_u0)
syncEnable_u361_u0<={add_u1132[31:4], 4'b10};
end
always @(posedge CLK)
begin
if (and_u2619_u0)
syncEnable_u362_u0<={add_u1136[31:4], 4'b10};
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_result_delayed_u7_u0<=1'h0;
else block_GO_delayed_result_delayed_u7_u0<=block_GO_delayed_u41_u0;
end
always @(posedge CLK)
begin
if (and_u2619_u0)
syncEnable_u363_u0<={add_u1128[31:4], 4'b1110};
end
always @(posedge CLK)
begin
if (and_u2619_u0)
syncEnable_u364_u0<={add_u1124[31:4], 4'b1110};
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01cf1df3_u0<=1'h0;
else reg_01cf1df3_u0<=and_delayed_result_delayed_u11_u0;
end
assign lessThanEqualTo_u11_a_signed=mux_u487_u0;
assign lessThanEqualTo_u11_b_signed=32'h37;
assign lessThanEqualTo_u11=lessThanEqualTo_u11_a_signed<=lessThanEqualTo_u11_b_signed;
assign not_u548_u0=~lessThanEqualTo_u11;
assign and_u2626_u0=or_u728_u0&lessThanEqualTo_u11;
assign and_u2627_u0=or_u728_u0&not_u548_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_u11_u0<=1'h0;
else and_delayed_result_delayed_u11_u0<=and_delayed_u63_u0;
end
assign and_u2628_u0=and_u2627_u0&or_u728_u0;
assign latch_01b87821_out=(and_u2618_u0)?32'h1e:32'h1e;
always @(posedge CLK)
begin
if (and_u2618_u0)
latch_01b87821_reg<=6'h1e;
end
assign latch_006cd68c_out=(and_u2618_u0)?32'h37:32'h37;
always @(posedge CLK)
begin
if (and_u2618_u0)
latch_006cd68c_reg<=7'h37;
end
assign mux_u487_u0=(reg_01cf1df3_u0)?syncEnable_u360_u0:32'h19;
assign latch_0083bde1_out=(and_u2618_u0)?32'h32:32'h32;
always @(posedge CLK)
begin
if (and_u2618_u0)
latch_0083bde1_reg<=7'h32;
end
assign or_u728_u0=reg_01cf1df3_u0|and_u2618_u0;
assign mux_u488_u0=(block_GO_delayed_result_delayed_u6)?syncEnable_u354_u0:{syncEnable_u361_u0[31:4], 4'b10};
assign or_u729_u0=block_GO_delayed_result_delayed_u6|block_GO_delayed_result_delayed_u7_u0;
assign or_u730_u0=block_GO_delayed_u40|block_GO_delayed_u41_u0;
assign mux_u489_u0=(block_GO_delayed_u40)?syncEnable_u355_u0:{syncEnable_u364_u0[31:4], 4'b1110};
assign or_u731_u0=block_GO_delayed_result_delayed_u6|block_GO_delayed_result_delayed_u7_u0;
assign mux_u490_u0=(block_GO_delayed_result_delayed_u6)?syncEnable_u352_u0:{syncEnable_u359_u0[31:4], 4'b10};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_017046c7_u0<=1'h0;
else reg_017046c7_u0<=GO;
end
assign mux_u491_u0=(block_GO_delayed_result_delayed_u6)?syncEnable_u356_u0:{syncEnable_u362_u0[31:4], 4'b10};
assign or_u732_u0=block_GO_delayed_result_delayed_u6|block_GO_delayed_result_delayed_u7_u0;
assign or_u733_u0=block_GO_delayed_u40|block_GO_delayed_u41_u0;
assign mux_u492_u0=(block_GO_delayed_u40)?syncEnable_u353_u0:{syncEnable_u363_u0[31:4], 4'b1110};
assign or_u734_u0=block_GO_delayed_u40|block_GO_delayed_u41_u0;
assign mux_u493_u0=(block_GO_delayed_u40)?syncEnable_u357_u0:{syncEnable_u358_u0[31:4], 4'b1110};
assign RESULT=or_u730_u0;
assign RESULT_u1914=mux_u489_u0;
assign RESULT_u1915=8'h0;
assign RESULT_u1916=3'h1;
assign RESULT_u1917=or_u733_u0;
assign RESULT_u1918=mux_u492_u0;
assign RESULT_u1919=8'h0;
assign RESULT_u1920=3'h1;
assign RESULT_u1921=or_u731_u0;
assign RESULT_u1922=mux_u490_u0;
assign RESULT_u1923=8'h0;
assign RESULT_u1924=3'h1;
assign RESULT_u1925=or_u734_u0;
assign RESULT_u1926=mux_u493_u0;
assign RESULT_u1927=8'hff;
assign RESULT_u1928=3'h1;
assign RESULT_u1929=or_u729_u0;
assign RESULT_u1930=mux_u488_u0;
assign RESULT_u1931=8'hff;
assign RESULT_u1932=3'h1;
assign RESULT_u1933=or_u732_u0;
assign RESULT_u1934=mux_u491_u0;
assign RESULT_u1935=8'h0;
assign RESULT_u1936=3'h1;
assign DONE=and_u2628_u0;
endmodule



module Generation_stateVar_state_s0(bus_0122c06d_, bus_00873bde_, bus_011920d6_, bus_0020f994_, bus_01530c78_);
input		bus_0122c06d_;
input		bus_00873bde_;
input		bus_011920d6_;
input		bus_0020f994_;
output		bus_01530c78_;
reg		stateVar_state_s0_u34=1'h0;
assign bus_01530c78_=stateVar_state_s0_u34;
always @(posedge bus_0122c06d_ or posedge bus_00873bde_)
begin
if (bus_00873bde_)
stateVar_state_s0_u34<=1'h0;
else if (bus_011920d6_)
stateVar_state_s0_u34<=bus_0020f994_;
end
endmodule



module Generation_getValueRGB(CLK, RESET, GO, port_007bdc5b_, port_01263d81_, port_01f1afae_, port_000d5d4f_, port_009075e0_, port_004cc74e_, port_0040ae5e_, port_00960a11_, RESULT, RESULT_u1937, RESULT_u1938, RESULT_u1939, RESULT_u1940, RESULT_u1941, RESULT_u1942, RESULT_u1943, RESULT_u1944, RESULT_u1945, RESULT_u1946, RESULT_u1947, RESULT_u1948, RESULT_u1949, RESULT_u1950, RESULT_u1951, RESULT_u1952, RESULT_u1953, RESULT_u1954, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_007bdc5b_;
input	[31:0]	port_01263d81_;
input		port_01f1afae_;
input		port_000d5d4f_;
input		port_009075e0_;
input	[7:0]	port_004cc74e_;
input	[7:0]	port_0040ae5e_;
input	[7:0]	port_00960a11_;
output		RESULT;
output	[31:0]	RESULT_u1937;
output		RESULT_u1938;
output	[31:0]	RESULT_u1939;
output		RESULT_u1940;
output	[31:0]	RESULT_u1941;
output	[7:0]	RESULT_u1942;
output	[2:0]	RESULT_u1943;
output		RESULT_u1944;
output	[31:0]	RESULT_u1945;
output	[7:0]	RESULT_u1946;
output	[2:0]	RESULT_u1947;
output		RESULT_u1948;
output	[31:0]	RESULT_u1949;
output	[7:0]	RESULT_u1950;
output	[2:0]	RESULT_u1951;
output		RESULT_u1952;
output		RESULT_u1953;
output		RESULT_u1954;
output		DONE;
wire		simplePinWrite;
wire		simplePinWrite_u700;
wire		simplePinWrite_u701;
wire	[31:0]	add;
wire	[31:0]	add_u1142;
wire	[31:0]	add_u1143;
wire	[31:0]	add_u1144;
wire		or_u735_u0;
reg		reg_01638321_u0=1'h0;
wire		and_u2629_u0;
wire	[31:0]	add_u1145;
wire	[31:0]	add_u1146;
wire	[31:0]	add_u1147;
wire	[31:0]	add_u1148;
wire		and_u2630_u0;
wire		or_u736_u0;
reg		reg_003dbe40_u0=1'h0;
wire	[31:0]	add_u1149;
wire	[31:0]	add_u1150;
wire	[31:0]	add_u1151;
wire	[31:0]	add_u1152;
reg		reg_01477fbb_u0=1'h0;
wire		or_u737_u0;
wire		and_u2631_u0;
wire	[31:0]	add_u1153;
wire signed	[31:0]	equals_b_signed;
wire		equals;
wire signed	[31:0]	equals_a_signed;
wire		and_u2632_u0;
wire		not_u549_u0;
wire		and_u2633_u0;
wire	[31:0]	add_u1154;
wire		and_u2634_u0;
wire	[31:0]	mux_u494;
wire	[31:0]	mux_u495_u0;
wire		and_u2635_u0;
reg	[31:0]	syncEnable_u365=32'h0;
reg	[7:0]	syncEnable_u366_u0=8'h0;
reg	[7:0]	syncEnable_u367_u0=8'h0;
reg		reg_0060a90c_u0=1'h0;
reg	[31:0]	syncEnable_u368_u0=32'h0;
reg	[31:0]	syncEnable_u369_u0=32'h0;
reg		reg_01b45de3_u0=1'h0;
reg	[7:0]	syncEnable_u370_u0=8'h0;
assign simplePinWrite=GO&{1{GO}};
assign simplePinWrite_u700=GO&{1{GO}};
assign simplePinWrite_u701=GO&{1{GO}};
assign add={port_007bdc5b_[24:0], 7'b0}+{port_007bdc5b_[26:0], 5'b0};
assign add_u1142={add[31:5], 5'b0}+{port_007bdc5b_[27:0], 4'b0};
assign add_u1143={add_u1142[31:4], 4'b0}+port_01263d81_;
assign add_u1144=32'h0+add_u1143;
assign or_u735_u0=and_u2629_u0|RESET;
always @(posedge CLK or posedge reg_01b45de3_u0 or posedge or_u735_u0)
begin
if (or_u735_u0)
reg_01638321_u0<=1'h0;
else if (reg_01b45de3_u0)
reg_01638321_u0<=1'h1;
else reg_01638321_u0<=reg_01638321_u0;
end
assign and_u2629_u0=reg_01638321_u0&port_009075e0_;
assign add_u1145={port_007bdc5b_[24:0], 7'b0}+{port_007bdc5b_[26:0], 5'b0};
assign add_u1146={add_u1145[31:5], 5'b0}+{port_007bdc5b_[27:0], 4'b0};
assign add_u1147={add_u1146[31:4], 4'b0}+port_01263d81_;
assign add_u1148=32'h0+add_u1147;
assign and_u2630_u0=reg_003dbe40_u0&port_000d5d4f_;
assign or_u736_u0=and_u2630_u0|RESET;
always @(posedge CLK or posedge reg_01b45de3_u0 or posedge or_u736_u0)
begin
if (or_u736_u0)
reg_003dbe40_u0<=1'h0;
else if (reg_01b45de3_u0)
reg_003dbe40_u0<=1'h1;
else reg_003dbe40_u0<=reg_003dbe40_u0;
end
assign add_u1149={port_007bdc5b_[24:0], 7'b0}+{port_007bdc5b_[26:0], 5'b0};
assign add_u1150={add_u1149[31:5], 5'b0}+{port_007bdc5b_[27:0], 4'b0};
assign add_u1151={add_u1150[31:4], 4'b0}+port_01263d81_;
assign add_u1152=32'h0+add_u1151;
always @(posedge CLK or posedge reg_01b45de3_u0 or posedge or_u737_u0)
begin
if (or_u737_u0)
reg_01477fbb_u0<=1'h0;
else if (reg_01b45de3_u0)
reg_01477fbb_u0<=1'h1;
else reg_01477fbb_u0<=reg_01477fbb_u0;
end
assign or_u737_u0=and_u2631_u0|RESET;
assign and_u2631_u0=reg_01477fbb_u0&port_01f1afae_;
assign add_u1153=port_01263d81_+32'h1;
assign equals_a_signed=add_u1153;
assign equals_b_signed=32'hb0;
assign equals=equals_a_signed==equals_b_signed;
assign and_u2632_u0=GO&not_u549_u0;
assign not_u549_u0=~equals;
assign and_u2633_u0=GO&equals;
assign add_u1154=port_007bdc5b_+32'h1;
assign and_u2634_u0=and_u2633_u0&GO;
assign mux_u494=(and_u2635_u0)?add_u1153:32'h0;
assign mux_u495_u0=(and_u2635_u0)?port_007bdc5b_:add_u1154;
assign and_u2635_u0=and_u2632_u0&GO;
always @(posedge CLK)
begin
if (GO)
syncEnable_u365<=add_u1152;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u366_u0<=port_00960a11_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u367_u0<=port_0040ae5e_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0060a90c_u0<=1'h0;
else reg_0060a90c_u0<=reg_01b45de3_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u368_u0<=add_u1144;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u369_u0<=add_u1148;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01b45de3_u0<=1'h0;
else reg_01b45de3_u0<=GO;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u370_u0<=port_004cc74e_;
end
assign RESULT=GO;
assign RESULT_u1937=mux_u495_u0;
assign RESULT_u1938=GO;
assign RESULT_u1939=mux_u494;
assign RESULT_u1940=reg_01b45de3_u0;
assign RESULT_u1941=syncEnable_u365;
assign RESULT_u1942=syncEnable_u367_u0;
assign RESULT_u1943=3'h1;
assign RESULT_u1944=reg_01b45de3_u0;
assign RESULT_u1945=syncEnable_u369_u0;
assign RESULT_u1946=syncEnable_u370_u0;
assign RESULT_u1947=3'h1;
assign RESULT_u1948=reg_01b45de3_u0;
assign RESULT_u1949=syncEnable_u368_u0;
assign RESULT_u1950=syncEnable_u366_u0;
assign RESULT_u1951=3'h1;
assign RESULT_u1952=simplePinWrite_u701;
assign RESULT_u1953=simplePinWrite;
assign RESULT_u1954=simplePinWrite_u700;
assign DONE=reg_0060a90c_u0;
endmodule



module Generation_Kicker_57(CLK, RESET, bus_00c4eeea_);
input		CLK;
input		RESET;
output		bus_00c4eeea_;
wire		bus_00070e49_;
reg		kicker_1=1'h0;
wire		bus_0173de00_;
wire		bus_00cef502_;
reg		kicker_2=1'h0;
reg		kicker_res=1'h0;
wire		bus_00e75e4e_;
assign bus_00070e49_=~RESET;
always @(posedge CLK)
begin
kicker_1<=bus_00070e49_;
end
assign bus_0173de00_=kicker_1&bus_00070e49_&bus_00e75e4e_;
assign bus_00cef502_=bus_00070e49_&kicker_1;
always @(posedge CLK)
begin
kicker_2<=bus_00cef502_;
end
always @(posedge CLK)
begin
kicker_res<=bus_0173de00_;
end
assign bus_00e75e4e_=~kicker_2;
assign bus_00c4eeea_=kicker_res;
endmodule



module Generation_stateVar_state_s2(bus_0168a69b_, bus_01920bdc_, bus_0105be8f_, bus_01b9532b_, bus_01ad823d_);
input		bus_0168a69b_;
input		bus_01920bdc_;
input		bus_0105be8f_;
input		bus_01b9532b_;
output		bus_01ad823d_;
reg		stateVar_state_s2_u32=1'h0;
assign bus_01ad823d_=stateVar_state_s2_u32;
always @(posedge bus_0168a69b_ or posedge bus_01920bdc_)
begin
if (bus_01920bdc_)
stateVar_state_s2_u32<=1'h0;
else if (bus_0105be8f_)
stateVar_state_s2_u32<=bus_01b9532b_;
end
endmodule



module Generation_forge_memory_25344x8_75(CLK, ENA, WEA, DINA, ENB, WEB, DINB, ADDRA, ADDRB, DOUTA, DONEA, DONEB);
input		CLK;
input		ENA;
input		WEA;
input	[7:0]	DINA;
input		ENB;
input		WEB;
input	[7:0]	DINB;
input	[31:0]	ADDRA;
input	[31:0]	ADDRB;
output	[7:0]	DOUTA;
output		DONEA;
output		DONEB;
wire		wea_0;
wire		web_0;
wire	[7:0]	pre_douta_0;
wire		wea_1;
wire		web_1;
wire	[7:0]	pre_douta_1;
reg	[7:0]	mux_outa;
reg	[31:0]	ADDRA_reg;
reg	[31:0]	ADDRB_reg;
wire	[7:0]	pre_doutb_1;
reg	[7:0]	mux_outb;
wire	[7:0]	pre_doutb_0;
reg		wea_done;
reg		rea_done;
reg		web_done;
assign wea_0=WEA&(ADDRA[31:14]==18'h0);
assign web_0=WEB&(ADDRB[31:14]==18'h0);
assign wea_1=WEA&(ADDRA[31:14]==18'h1);
assign web_1=WEB&(ADDRB[31:14]==18'h1);
always @(posedge CLK)
begin
ADDRA_reg<=ADDRA;
end
always @(ADDRA_reg or pre_douta_0 or pre_douta_1)
begin
case (ADDRA_reg[31:14])18'd0:mux_outa=pre_douta_0;
18'd1:mux_outa=pre_douta_1;
default:mux_outa=8'h0;
endcase end
always @(posedge CLK)
begin
ADDRB_reg<=ADDRB;
end
always @(ADDRB_reg or pre_doutb_0 or pre_doutb_1)
begin
case (ADDRB_reg[31:14])18'd0:mux_outb=pre_doutb_0;
18'd1:mux_outb=pre_doutb_1;
default:mux_outb=8'h0;
endcase end
always @(posedge CLK)
begin
wea_done<=WEA;
rea_done<=ENA;
web_done<=WEB;
end
assign DONEA=wea_done|rea_done;
assign DONEB=web_done;
assign DOUTA=mux_outa;
// Memory array element: COL: 0, ROW: 0
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_272(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[0]), .DOA(pre_douta_0[0]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[0]), .DOB());
// Memory array element: COL: 0, ROW: 1
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_273(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[1]), .DOA(pre_douta_0[1]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[1]), .DOB());
// Memory array element: COL: 0, ROW: 2
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_274(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[2]), .DOA(pre_douta_0[2]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[2]), .DOB());
// Memory array element: COL: 0, ROW: 3
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_275(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[3]), .DOA(pre_douta_0[3]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[3]), .DOB());
// Memory array element: COL: 0, ROW: 4
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_276(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[4]), .DOA(pre_douta_0[4]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[4]), .DOB());
// Memory array element: COL: 0, ROW: 5
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_277(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[5]), .DOA(pre_douta_0[5]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[5]), .DOB());
// Memory array element: COL: 0, ROW: 6
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_278(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[6]), .DOA(pre_douta_0[6]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[6]), .DOB());
// Memory array element: COL: 0, ROW: 7
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_279(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[7]), .DOA(pre_douta_0[7]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[7]), .DOB());
// Memory array element: COL: 1, ROW: 0
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_280(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[0]), .DOA(pre_douta_1[0]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[0]), .DOB());
// Memory array element: COL: 1, ROW: 1
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_281(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[1]), .DOA(pre_douta_1[1]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[1]), .DOB());
// Memory array element: COL: 1, ROW: 2
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_282(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[2]), .DOA(pre_douta_1[2]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[2]), .DOB());
// Memory array element: COL: 1, ROW: 3
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_283(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[3]), .DOA(pre_douta_1[3]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[3]), .DOB());
// Memory array element: COL: 1, ROW: 4
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_284(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[4]), .DOA(pre_douta_1[4]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[4]), .DOB());
// Memory array element: COL: 1, ROW: 5
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_285(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[5]), .DOA(pre_douta_1[5]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[5]), .DOB());
// Memory array element: COL: 1, ROW: 6
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_286(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[6]), .DOA(pre_douta_1[6]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[6]), .DOB());
// Memory array element: COL: 1, ROW: 7
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_287(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[7]), .DOA(pre_douta_1[7]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[7]), .DOB());
endmodule



module Generation_structuralmemory_0156af01_(CLK_u49, bus_0073ced7_, bus_00fc033f_, bus_00b8b050_, bus_0140811d_, bus_008c32f9_, bus_002bf4e6_, bus_00a404ce_, bus_0192694e_, bus_0141e826_, bus_00d571fa_, bus_01dc999c_, bus_01db46e6_, bus_012df243_);
input		CLK_u49;
input		bus_0073ced7_;
input	[31:0]	bus_00fc033f_;
input	[2:0]	bus_00b8b050_;
input		bus_0140811d_;
input		bus_008c32f9_;
input	[7:0]	bus_002bf4e6_;
input	[31:0]	bus_00a404ce_;
input	[2:0]	bus_0192694e_;
input		bus_0141e826_;
input	[7:0]	bus_00d571fa_;
output	[7:0]	bus_01dc999c_;
output		bus_01db46e6_;
output		bus_012df243_;
wire		or_012bb3fe_u0;
reg		logicalMem_159414f_re_delay0_u0=1'h0;
reg		logicalMem_159414f_we_delay0_u0=1'h0;
reg		logicalMem_159414f_we_delay0_u1_u0=1'h0;
wire	[7:0]	bus_01ccde21_;
wire		or_015fa1fb_u0;
assign or_012bb3fe_u0=logicalMem_159414f_re_delay0_u0|logicalMem_159414f_we_delay0_u0;
assign bus_01dc999c_=bus_01ccde21_;
assign bus_01db46e6_=or_012bb3fe_u0;
assign bus_012df243_=logicalMem_159414f_we_delay0_u1_u0;
always @(posedge CLK_u49 or posedge bus_0073ced7_)
begin
if (bus_0073ced7_)
logicalMem_159414f_re_delay0_u0<=1'h0;
else logicalMem_159414f_re_delay0_u0<=bus_0140811d_;
end
always @(posedge CLK_u49 or posedge bus_0073ced7_)
begin
if (bus_0073ced7_)
logicalMem_159414f_we_delay0_u0<=1'h0;
else logicalMem_159414f_we_delay0_u0<=bus_008c32f9_;
end
always @(posedge CLK_u49 or posedge bus_0073ced7_)
begin
if (bus_0073ced7_)
logicalMem_159414f_we_delay0_u1_u0<=1'h0;
else logicalMem_159414f_we_delay0_u1_u0<=bus_0141e826_;
end
Generation_forge_memory_25344x8_75 Generation_forge_memory_25344x8_75_instance0(.CLK(CLK_u49), 
  .ENA(or_015fa1fb_u0), .WEA(bus_008c32f9_), .DINA(bus_002bf4e6_), .ADDRA(bus_00fc033f_), 
  .DOUTA(bus_01ccde21_), .DONEA(), .ENB(bus_0141e826_), .WEB(bus_0141e826_), .DINB(8'hff), 
  .ADDRB(bus_00a404ce_), .DONEB());
assign or_015fa1fb_u0=bus_0140811d_|bus_008c32f9_;
endmodule



module Generation_doneCountIm(CLK, RESET, GO, RESULT, RESULT_u1955, DONE);
input		CLK;
input		RESET;
input		GO;
output		RESULT;
output	[31:0]	RESULT_u1955;
output		DONE;
reg		reg_0094d112_u0=1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0094d112_u0<=1'h0;
else reg_0094d112_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u1955=32'h0;
assign DONE=reg_0094d112_u0;
endmodule



module Generation_simplememoryreferee_000742eb_(bus_0019d89f_, bus_00dcc243_, bus_0057a34a_, bus_013da532_, bus_00660791_, bus_007fe65e_, bus_01d1ac5f_, bus_01679577_, bus_00287f7c_, bus_01867765_, bus_0136da55_, bus_0086d7cf_, bus_01fe6336_, bus_0185bd7a_);
input		bus_0019d89f_;
input		bus_00dcc243_;
input		bus_0057a34a_;
input	[7:0]	bus_013da532_;
input		bus_00660791_;
input	[7:0]	bus_007fe65e_;
input	[31:0]	bus_01d1ac5f_;
input	[2:0]	bus_01679577_;
output	[7:0]	bus_00287f7c_;
output	[31:0]	bus_01867765_;
output		bus_0136da55_;
output		bus_0086d7cf_;
output	[2:0]	bus_01fe6336_;
output		bus_0185bd7a_;
assign bus_00287f7c_=8'h0;
assign bus_01867765_=bus_01d1ac5f_;
assign bus_0136da55_=bus_00660791_;
assign bus_0086d7cf_=bus_00660791_;
assign bus_01fe6336_=3'h1;
assign bus_0185bd7a_=bus_0057a34a_;
endmodule



module Generation_structuralmemory_00c0d3f6_(CLK_u50, bus_01d2754e_, bus_000dbf39_, bus_0149775b_, bus_003a8ec4_, bus_01674500_, bus_0108036b_, bus_01ae55ef_, bus_00a5d728_, bus_01563c6d_, bus_000f6b16_, bus_0072ed28_, bus_01188a3b_, bus_003f9e84_);
input		CLK_u50;
input		bus_01d2754e_;
input	[31:0]	bus_000dbf39_;
input	[2:0]	bus_0149775b_;
input		bus_003a8ec4_;
input		bus_01674500_;
input	[7:0]	bus_0108036b_;
input	[31:0]	bus_01ae55ef_;
input	[2:0]	bus_00a5d728_;
input		bus_01563c6d_;
input	[7:0]	bus_000f6b16_;
output	[7:0]	bus_0072ed28_;
output		bus_01188a3b_;
output		bus_003f9e84_;
reg		logicalMem_e7beaf_we_delay0_u0=1'h0;
wire		or_01bb871f_u0;
wire		or_01fda1b9_u0;
reg		logicalMem_e7beaf_re_delay0_u0=1'h0;
wire	[7:0]	bus_01876f43_;
reg		logicalMem_e7beaf_we_delay0_u1_u0=1'h0;
always @(posedge CLK_u50 or posedge bus_01d2754e_)
begin
if (bus_01d2754e_)
logicalMem_e7beaf_we_delay0_u0<=1'h0;
else logicalMem_e7beaf_we_delay0_u0<=bus_01674500_;
end
assign bus_0072ed28_=bus_01876f43_;
assign bus_01188a3b_=or_01fda1b9_u0;
assign bus_003f9e84_=logicalMem_e7beaf_we_delay0_u1_u0;
assign or_01bb871f_u0=bus_003a8ec4_|bus_01674500_;
assign or_01fda1b9_u0=logicalMem_e7beaf_re_delay0_u0|logicalMem_e7beaf_we_delay0_u0;
always @(posedge CLK_u50 or posedge bus_01d2754e_)
begin
if (bus_01d2754e_)
logicalMem_e7beaf_re_delay0_u0<=1'h0;
else logicalMem_e7beaf_re_delay0_u0<=bus_003a8ec4_;
end
Generation_forge_memory_25344x8_75 Generation_forge_memory_25344x8_75_instance1(.CLK(CLK_u50), 
  .ENA(or_01bb871f_u0), .WEA(bus_01674500_), .DINA(bus_0108036b_), .ADDRA(bus_000dbf39_), 
  .DOUTA(bus_01876f43_), .DONEA(), .ENB(bus_01563c6d_), .WEB(bus_01563c6d_), .DINB(8'h0), 
  .ADDRB(bus_01ae55ef_), .DONEB());
always @(posedge CLK_u50 or posedge bus_01d2754e_)
begin
if (bus_01d2754e_)
logicalMem_e7beaf_we_delay0_u1_u0<=1'h0;
else logicalMem_e7beaf_we_delay0_u1_u0<=bus_01563c6d_;
end
endmodule



module Generation_globalreset_physical_018187f8_(bus_00cbf5a7_, bus_0058fdd8_, bus_01d34608_);
input		bus_00cbf5a7_;
input		bus_0058fdd8_;
output		bus_01d34608_;
reg		glitch_u57=1'h0;
wire		and_017eccba_u0;
wire		or_0081a152_u0;
wire		not_00c85999_u0;
reg		final_u57=1'h1;
reg		cross_u57=1'h0;
reg		sample_u57=1'h0;
always @(posedge bus_00cbf5a7_)
begin
glitch_u57<=cross_u57;
end
assign and_017eccba_u0=cross_u57&glitch_u57;
assign bus_01d34608_=or_0081a152_u0;
assign or_0081a152_u0=bus_0058fdd8_|final_u57;
assign not_00c85999_u0=~and_017eccba_u0;
always @(posedge bus_00cbf5a7_)
begin
final_u57<=not_00c85999_u0;
end
always @(posedge bus_00cbf5a7_)
begin
cross_u57<=sample_u57;
end
always @(posedge bus_00cbf5a7_)
begin
sample_u57<=1'h1;
end
endmodule



module Generation_simplememoryreferee_0062bad9_(bus_006120d5_, bus_00b2b57c_, bus_018943bd_, bus_007f922a_, bus_0128b244_, bus_01da6bec_, bus_00a675df_, bus_00b36d07_, bus_011ac12c_, bus_004c87c7_, bus_01fc3728_, bus_005db036_, bus_01966503_, bus_005f1004_, bus_00837cdf_, bus_015536f1_, bus_004d0152_, bus_01d90de5_, bus_0042f76c_, bus_015b9c7d_, bus_01bb2165_, bus_00dbd379_, bus_00c1d8fc_, bus_007b17d0_);
input		bus_006120d5_;
input		bus_00b2b57c_;
input		bus_018943bd_;
input	[7:0]	bus_007f922a_;
input		bus_0128b244_;
input	[7:0]	bus_01da6bec_;
input	[31:0]	bus_00a675df_;
input	[2:0]	bus_00b36d07_;
input		bus_011ac12c_;
input	[7:0]	bus_004c87c7_;
input	[31:0]	bus_01fc3728_;
input	[2:0]	bus_005db036_;
input		bus_01966503_;
input	[31:0]	bus_005f1004_;
input	[2:0]	bus_00837cdf_;
output	[7:0]	bus_015536f1_;
output	[31:0]	bus_004d0152_;
output		bus_01d90de5_;
output		bus_0042f76c_;
output	[2:0]	bus_015b9c7d_;
output		bus_01bb2165_;
output		bus_00dbd379_;
output	[7:0]	bus_00c1d8fc_;
output		bus_007b17d0_;
reg		done_qual_u150_u0=1'h0;
wire		not_0107ee33_u0;
reg		done_qual_u151_u0=1'h0;
wire		or_00a3edc2_u0;
wire		or_01ec1c11_u0;
wire		or_0137dfd5_u0;
wire		and_01699b24_u0;
wire		not_01e13dba_u0;
wire		or_0034a7e6_u0;
wire		and_00cd0836_u0;
wire	[31:0]	mux_0053f438_u0;
wire		and_00daf273_u0;
reg		done_qual_u152_u0=1'h0;
wire		or_01e56e51_u0;
wire		not_01b51865_u0;
wire	[7:0]	mux_01afa376_u0;
always @(posedge bus_006120d5_)
begin
if (bus_00b2b57c_)
done_qual_u150_u0<=1'h0;
else done_qual_u150_u0<=bus_01966503_;
end
assign not_0107ee33_u0=~bus_018943bd_;
always @(posedge bus_006120d5_)
begin
if (bus_00b2b57c_)
done_qual_u151_u0<=1'h0;
else done_qual_u151_u0<=bus_0128b244_;
end
assign or_00a3edc2_u0=bus_011ac12c_|done_qual_u152_u0;
assign or_01ec1c11_u0=bus_0128b244_|done_qual_u151_u0;
assign or_0137dfd5_u0=bus_01966503_|done_qual_u150_u0;
assign and_01699b24_u0=or_00a3edc2_u0&bus_018943bd_;
assign not_01e13dba_u0=~bus_018943bd_;
assign or_0034a7e6_u0=bus_0128b244_|bus_011ac12c_;
assign and_00cd0836_u0=or_01ec1c11_u0&bus_018943bd_;
assign mux_0053f438_u0=({32{bus_0128b244_}}&bus_00a675df_)|({32{bus_011ac12c_}}&bus_01fc3728_)|({32{bus_01966503_}}&bus_005f1004_);
assign and_00daf273_u0=or_0137dfd5_u0&bus_018943bd_;
always @(posedge bus_006120d5_)
begin
if (bus_00b2b57c_)
done_qual_u152_u0<=1'h0;
else done_qual_u152_u0<=bus_011ac12c_;
end
assign or_01e56e51_u0=bus_0128b244_|bus_011ac12c_|bus_01966503_;
assign not_01b51865_u0=~bus_018943bd_;
assign mux_01afa376_u0=(bus_0128b244_)?bus_01da6bec_:8'h0;
assign bus_015536f1_=mux_01afa376_u0;
assign bus_004d0152_=mux_0053f438_u0;
assign bus_01d90de5_=or_0034a7e6_u0;
assign bus_0042f76c_=or_01e56e51_u0;
assign bus_015b9c7d_=3'h1;
assign bus_01bb2165_=and_00cd0836_u0;
assign bus_00dbd379_=and_01699b24_u0;
assign bus_00c1d8fc_=bus_007f922a_;
assign bus_007b17d0_=and_00daf273_u0;
endmodule



module Generation_endianswapper_0024d79b_(endianswapper_0024d79b_in, endianswapper_0024d79b_out);
input	[31:0]	endianswapper_0024d79b_in;
output	[31:0]	endianswapper_0024d79b_out;
assign endianswapper_0024d79b_out=endianswapper_0024d79b_in;
endmodule



module Generation_endianswapper_01d49a44_(endianswapper_01d49a44_in, endianswapper_01d49a44_out);
input	[31:0]	endianswapper_01d49a44_in;
output	[31:0]	endianswapper_01d49a44_out;
assign endianswapper_01d49a44_out=endianswapper_01d49a44_in;
endmodule



module Generation_stateVar_count_y(bus_0168294f_, bus_017039a6_, bus_0130359b_, bus_00d547ca_, bus_007d4ec1_, bus_00272892_, bus_00e65a1a_);
input		bus_0168294f_;
input		bus_017039a6_;
input		bus_0130359b_;
input	[31:0]	bus_00d547ca_;
input		bus_007d4ec1_;
input	[31:0]	bus_00272892_;
output	[31:0]	bus_00e65a1a_;
wire		or_01d9785c_u0;
wire	[31:0]	endianswapper_0024d79b_out;
reg	[31:0]	stateVar_count_y_u11=32'h0;
wire	[31:0]	mux_01300c66_u0;
wire	[31:0]	endianswapper_01d49a44_out;
assign or_01d9785c_u0=bus_0130359b_|bus_007d4ec1_;
Generation_endianswapper_0024d79b_ Generation_endianswapper_0024d79b__1(.endianswapper_0024d79b_in(stateVar_count_y_u11), 
  .endianswapper_0024d79b_out(endianswapper_0024d79b_out));
always @(posedge bus_0168294f_ or posedge bus_017039a6_)
begin
if (bus_017039a6_)
stateVar_count_y_u11<=32'h0;
else if (or_01d9785c_u0)
stateVar_count_y_u11<=endianswapper_01d49a44_out;
end
assign bus_00e65a1a_=endianswapper_0024d79b_out;
assign mux_01300c66_u0=(bus_0130359b_)?bus_00d547ca_:bus_00272892_;
Generation_endianswapper_01d49a44_ Generation_endianswapper_01d49a44__1(.endianswapper_01d49a44_in(mux_01300c66_u0), 
  .endianswapper_01d49a44_out(endianswapper_01d49a44_out));
endmodule



module Generation_simplememoryreferee_01801ae8_(bus_005cefdf_, bus_01883661_, bus_01533ec6_, bus_01625b66_, bus_005222c2_, bus_004e4c93_, bus_008195d8_, bus_0133852a_, bus_005e8953_, bus_01465e99_, bus_01bd7297_, bus_0106a06d_, bus_005bc28e_, bus_016bc16f_);
input		bus_005cefdf_;
input		bus_01883661_;
input		bus_01533ec6_;
input	[7:0]	bus_01625b66_;
input		bus_005222c2_;
input	[7:0]	bus_004e4c93_;
input	[31:0]	bus_008195d8_;
input	[2:0]	bus_0133852a_;
output	[7:0]	bus_005e8953_;
output	[31:0]	bus_01465e99_;
output		bus_01bd7297_;
output		bus_0106a06d_;
output	[2:0]	bus_005bc28e_;
output		bus_016bc16f_;
assign bus_005e8953_=8'h0;
assign bus_01465e99_=bus_008195d8_;
assign bus_01bd7297_=bus_005222c2_;
assign bus_0106a06d_=bus_005222c2_;
assign bus_005bc28e_=3'h1;
assign bus_016bc16f_=bus_01533ec6_;
endmodule



module Generation_structuralmemory_01173ea4_(CLK_u51, bus_00145df3_, bus_012e52ce_, bus_0040491c_, bus_005d0e89_, bus_0041c93d_, bus_00133706_, bus_0085d248_, bus_00aaeacd_, bus_01b5bcf2_, bus_00bb37ab_, bus_016572b8_, bus_01818ac0_, bus_0143eb1d_);
input		CLK_u51;
input		bus_00145df3_;
input	[31:0]	bus_012e52ce_;
input	[2:0]	bus_0040491c_;
input		bus_005d0e89_;
input		bus_0041c93d_;
input	[7:0]	bus_00133706_;
input	[31:0]	bus_0085d248_;
input	[2:0]	bus_00aaeacd_;
input		bus_01b5bcf2_;
input	[7:0]	bus_00bb37ab_;
output	[7:0]	bus_016572b8_;
output		bus_01818ac0_;
output		bus_0143eb1d_;
reg		logicalMem_11fd73a_we_delay0_u0=1'h0;
wire		or_004777bf_u0;
reg		logicalMem_11fd73a_we_delay0_u1_u0=1'h0;
reg		logicalMem_11fd73a_re_delay0_u0=1'h0;
wire		or_00a12101_u0;
wire	[7:0]	bus_0195d60c_;
always @(posedge CLK_u51 or posedge bus_00145df3_)
begin
if (bus_00145df3_)
logicalMem_11fd73a_we_delay0_u0<=1'h0;
else logicalMem_11fd73a_we_delay0_u0<=bus_01b5bcf2_;
end
assign or_004777bf_u0=bus_005d0e89_|bus_0041c93d_;
assign bus_016572b8_=bus_0195d60c_;
assign bus_01818ac0_=or_00a12101_u0;
assign bus_0143eb1d_=logicalMem_11fd73a_we_delay0_u0;
always @(posedge CLK_u51 or posedge bus_00145df3_)
begin
if (bus_00145df3_)
logicalMem_11fd73a_we_delay0_u1_u0<=1'h0;
else logicalMem_11fd73a_we_delay0_u1_u0<=bus_0041c93d_;
end
always @(posedge CLK_u51 or posedge bus_00145df3_)
begin
if (bus_00145df3_)
logicalMem_11fd73a_re_delay0_u0<=1'h0;
else logicalMem_11fd73a_re_delay0_u0<=bus_005d0e89_;
end
assign or_00a12101_u0=logicalMem_11fd73a_re_delay0_u0|logicalMem_11fd73a_we_delay0_u1_u0;
Generation_forge_memory_25344x8_75 Generation_forge_memory_25344x8_75_instance2(.CLK(CLK_u51), 
  .ENA(or_004777bf_u0), .WEA(bus_0041c93d_), .DINA(bus_00133706_), .ADDRA(bus_012e52ce_), 
  .DOUTA(bus_0195d60c_), .DONEA(), .ENB(bus_01b5bcf2_), .WEB(bus_01b5bcf2_), .DINB(8'h0), 
  .ADDRB(bus_0085d248_), .DONEB());
endmodule



module Generation_simplememoryreferee_0173d745_(bus_00527630_, bus_01cd82ec_, bus_01248bfe_, bus_005611d2_, bus_00769b40_, bus_0149134b_, bus_0149fcb3_, bus_0148efea_, bus_0018bf4d_, bus_006f81ca_, bus_014b9e03_, bus_0065e7ab_, bus_00309326_, bus_01835b38_, bus_01b43d37_, bus_00ac07b4_, bus_00098098_, bus_003255c0_, bus_019964a1_, bus_00e47af6_, bus_017f06fa_, bus_004cb6d6_, bus_010ccceb_, bus_001efe58_);
input		bus_00527630_;
input		bus_01cd82ec_;
input		bus_01248bfe_;
input	[7:0]	bus_005611d2_;
input		bus_00769b40_;
input	[7:0]	bus_0149134b_;
input	[31:0]	bus_0149fcb3_;
input	[2:0]	bus_0148efea_;
input		bus_0018bf4d_;
input	[7:0]	bus_006f81ca_;
input	[31:0]	bus_014b9e03_;
input	[2:0]	bus_0065e7ab_;
input		bus_00309326_;
input	[31:0]	bus_01835b38_;
input	[2:0]	bus_01b43d37_;
output	[7:0]	bus_00ac07b4_;
output	[31:0]	bus_00098098_;
output		bus_003255c0_;
output		bus_019964a1_;
output	[2:0]	bus_00e47af6_;
output		bus_017f06fa_;
output		bus_004cb6d6_;
output	[7:0]	bus_010ccceb_;
output		bus_001efe58_;
wire		or_00564b7d_u0;
wire	[7:0]	mux_014579a3_u0;
wire		or_01ab2db1_u0;
reg		done_qual_u153_u0=1'h0;
reg		done_qual_u154_u0=1'h0;
wire		not_018d4523_u0;
wire		and_0023c09c_u0;
wire	[31:0]	mux_0174d087_u0;
wire		and_002245a0_u0;
wire		not_01f7bc60_u0;
wire		or_0010afa8_u0;
wire		or_01785a60_u0;
wire		or_001a7ade_u0;
reg		done_qual_u155_u0=1'h0;
wire		and_007f191e_u0;
wire		not_016804ac_u0;
assign or_00564b7d_u0=bus_00769b40_|bus_0018bf4d_;
assign mux_014579a3_u0=(bus_00769b40_)?bus_0149134b_:8'hff;
assign or_01ab2db1_u0=bus_00769b40_|done_qual_u154_u0;
always @(posedge bus_00527630_)
begin
if (bus_01cd82ec_)
done_qual_u153_u0<=1'h0;
else done_qual_u153_u0<=bus_0018bf4d_;
end
always @(posedge bus_00527630_)
begin
if (bus_01cd82ec_)
done_qual_u154_u0<=1'h0;
else done_qual_u154_u0<=bus_00769b40_;
end
assign not_018d4523_u0=~bus_01248bfe_;
assign and_0023c09c_u0=or_01ab2db1_u0&bus_01248bfe_;
assign mux_0174d087_u0=({32{bus_00769b40_}}&bus_0149fcb3_)|({32{bus_0018bf4d_}}&bus_014b9e03_)|({32{bus_00309326_}}&bus_01835b38_);
assign and_002245a0_u0=or_001a7ade_u0&bus_01248bfe_;
assign not_01f7bc60_u0=~bus_01248bfe_;
assign or_0010afa8_u0=bus_00769b40_|bus_0018bf4d_|bus_00309326_;
assign or_01785a60_u0=bus_00309326_|done_qual_u155_u0;
assign or_001a7ade_u0=bus_0018bf4d_|done_qual_u153_u0;
always @(posedge bus_00527630_)
begin
if (bus_01cd82ec_)
done_qual_u155_u0<=1'h0;
else done_qual_u155_u0<=bus_00309326_;
end
assign and_007f191e_u0=or_01785a60_u0&bus_01248bfe_;
assign bus_00ac07b4_=mux_014579a3_u0;
assign bus_00098098_=mux_0174d087_u0;
assign bus_003255c0_=or_00564b7d_u0;
assign bus_019964a1_=or_0010afa8_u0;
assign bus_00e47af6_=3'h1;
assign bus_017f06fa_=and_0023c09c_u0;
assign bus_004cb6d6_=and_002245a0_u0;
assign bus_010ccceb_=bus_005611d2_;
assign bus_001efe58_=and_007f191e_u0;
assign not_016804ac_u0=~bus_01248bfe_;
endmodule



module Generation_simplememoryreferee_00377ebe_(bus_014779db_, bus_01911ea6_, bus_019e8d0b_, bus_00efbc69_, bus_004c6569_, bus_007ef2a5_, bus_00d7d56a_, bus_0033b983_, bus_013a971b_, bus_011fbfd3_, bus_015957dd_, bus_0159ecfe_, bus_016e703b_, bus_01d84fc4_);
input		bus_014779db_;
input		bus_01911ea6_;
input		bus_019e8d0b_;
input	[7:0]	bus_00efbc69_;
input		bus_004c6569_;
input	[7:0]	bus_007ef2a5_;
input	[31:0]	bus_00d7d56a_;
input	[2:0]	bus_0033b983_;
output	[7:0]	bus_013a971b_;
output	[31:0]	bus_011fbfd3_;
output		bus_015957dd_;
output		bus_0159ecfe_;
output	[2:0]	bus_016e703b_;
output		bus_01d84fc4_;
assign bus_013a971b_=8'hff;
assign bus_011fbfd3_=bus_00d7d56a_;
assign bus_015957dd_=bus_004c6569_;
assign bus_0159ecfe_=bus_004c6569_;
assign bus_016e703b_=3'h1;
assign bus_01d84fc4_=bus_019e8d0b_;
endmodule



module Generation_scheduler(CLK, RESET, GO, port_0032333f_, port_01ce98f6_, port_00c47705_, port_00dad65c_, port_00a666cf_, port_012c5997_, port_001c856e_, port_000be277_, port_012fe075_, port_00d4319a_, port_00429cca_, port_00c133f5_, port_01d1c7ea_, port_010c32d0_, RESULT, RESULT_u1956, RESULT_u1957, RESULT_u1958, RESULT_u1959, RESULT_u1960, RESULT_u1961, RESULT_u1962, RESULT_u1963, RESULT_u1964, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_0032333f_;
input		port_01ce98f6_;
input		port_00c47705_;
input	[31:0]	port_00dad65c_;
input		port_00a666cf_;
input		port_012c5997_;
input		port_001c856e_;
input		port_000be277_;
input		port_012fe075_;
input		port_00d4319a_;
input		port_00429cca_;
input		port_00c133f5_;
input		port_01d1c7ea_;
input		port_010c32d0_;
output		RESULT;
output		RESULT_u1956;
output		RESULT_u1957;
output		RESULT_u1958;
output		RESULT_u1959;
output		RESULT_u1960;
output		RESULT_u1961;
output		RESULT_u1962;
output		RESULT_u1963;
output		RESULT_u1964;
output		DONE;
wire		and_u2636_u0;
wire		and_u2637_u0;
wire		and_u2638_u0;
wire		equals;
wire signed	[31:0]	equals_a_signed;
wire signed	[31:0]	equals_b_signed;
wire		and_u2639_u0;
wire		and_u2640_u0;
wire		not_u550_u0;
wire		and_u2641_u0;
wire		and_u2642_u0;
wire		and_u2643_u0;
wire		and_u2644_u0;
wire		not_u551_u0;
wire		simplePinWrite;
wire		and_u2645_u0;
wire		not_u552_u0;
wire		and_u2646_u0;
wire		and_u2647_u0;
wire		simplePinWrite_u702;
wire		and_u2648_u0;
reg		reg_002c1537_u0=1'h0;
wire		and_u2649_u0;
reg		reg_00ee82d4_u0=1'h0;
wire		or_u738_u0;
wire		and_u2650_u0;
reg		and_delayed_u64=1'h0;
wire		or_u739_u0;
reg		reg_00d4e6ed_u0=1'h0;
wire		and_u2651_u0;
wire		and_u2652_u0;
wire		or_u740_u0;
wire		and_u2653_u0;
reg		and_delayed_u65_u0=1'h0;
wire		and_u2654_u0;
wire		and_u2655_u0;
wire		not_u553_u0;
wire		and_u2656_u0;
wire		simplePinWrite_u703;
wire		and_u2657_u0;
wire		and_u2658_u0;
wire		or_u741_u0;
wire		and_u2659_u0;
reg		reg_00e338d7_u0=1'h0;
wire		and_u2660_u0;
wire		not_u554_u0;
wire		and_u2661_u0;
wire		and_u2662_u0;
wire		not_u555_u0;
wire		and_u2663_u0;
wire		and_u2664_u0;
wire		simplePinWrite_u704;
wire		and_u2665_u0;
wire		and_u2666_u0;
wire		and_u2667_u0;
wire		not_u556_u0;
wire		simplePinWrite_u705;
reg		reg_00cc41c6_u0=1'h0;
wire		or_u742_u0;
wire		and_u2668_u0;
reg		reg_001f57d1_u0=1'h0;
reg		reg_01d1ae03_u0=1'h0;
wire		and_u2669_u0;
wire		and_u2670_u0;
reg		reg_00f575f7_u0=1'h0;
wire		or_u743_u0;
wire		and_u2671_u0;
wire		and_u2672_u0;
wire		and_u2673_u0;
wire		and_u2674_u0;
wire		or_u744_u0;
reg		and_delayed_u66_u0=1'h0;
wire		mux_u496;
wire		or_u745_u0;
wire		mux_u497_u0;
wire		or_u746_u0;
wire		doneCountIm_go_merge;
wire		mux_u498_u0;
wire		or_u747_u0;
wire		scoreboard_00861902_resOr1;
wire		scoreboard_00861902_resOr0;
wire		bus_01994ea2_;
reg		scoreboard_00861902_reg0=1'h0;
reg		scoreboard_00861902_reg2=1'h0;
reg		scoreboard_00861902_reg1=1'h0;
wire		scoreboard_00861902_resOr2;
wire		scoreboard_00861902_and;
reg		syncEnable_u371=1'h0;
reg		syncEnable_u372_u0=1'h0;
reg		syncEnable_u373_u0=1'h0;
reg		block_GO_delayed_u42=1'h0;
reg		syncEnable_u374_u0=1'h0;
reg		syncEnable_u375_u0=1'h0;
wire		or_u748_u0;
reg		reg_0163200b_u0=1'h0;
wire		mux_u499_u0;
wire		or_u749_u0;
wire		mux_u500_u0;
wire		or_u750_u0;
reg		reg_0037d9b9_u0=1'h0;
wire		or_u751_u0;
wire		mux_u501_u0;
assign and_u2636_u0=or_u748_u0&or_u748_u0;
assign and_u2637_u0=port_00a666cf_&port_00c133f5_;
assign and_u2638_u0=and_u2637_u0&port_01d1c7ea_;
assign equals_a_signed=port_00dad65c_;
assign equals_b_signed=32'h90;
assign equals=equals_a_signed==equals_b_signed;
assign and_u2639_u0=port_001c856e_&port_000be277_;
assign and_u2640_u0=and_u2639_u0&port_00d4319a_;
assign not_u550_u0=~syncEnable_u372_u0;
assign and_u2641_u0=block_GO_delayed_u42&syncEnable_u372_u0;
assign and_u2642_u0=block_GO_delayed_u42&not_u550_u0;
assign and_u2643_u0=and_u2654_u0&not_u551_u0;
assign and_u2644_u0=and_u2654_u0&syncEnable_u371;
assign not_u551_u0=~syncEnable_u371;
assign simplePinWrite=and_u2645_u0&{1{and_u2645_u0}};
assign and_u2645_u0=and_u2651_u0&and_u2651_u0;
assign not_u552_u0=~syncEnable_u375_u0;
assign and_u2646_u0=and_u2652_u0&syncEnable_u375_u0;
assign and_u2647_u0=and_u2652_u0&not_u552_u0;
assign simplePinWrite_u702=and_u2648_u0&{1{and_u2648_u0}};
assign and_u2648_u0=and_u2649_u0&and_u2649_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_002c1537_u0<=1'h0;
else reg_002c1537_u0<=and_u2650_u0;
end
assign and_u2649_u0=and_u2646_u0&and_u2652_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00ee82d4_u0<=1'h0;
else reg_00ee82d4_u0<=and_delayed_u64;
end
assign or_u738_u0=reg_002c1537_u0|reg_00ee82d4_u0;
assign and_u2650_u0=and_u2647_u0&and_u2652_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u64<=1'h0;
else and_delayed_u64<=and_u2649_u0;
end
assign or_u739_u0=reg_00d4e6ed_u0|or_u738_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00d4e6ed_u0<=1'h0;
else reg_00d4e6ed_u0<=and_u2651_u0;
end
assign and_u2651_u0=and_u2644_u0&and_u2654_u0;
assign and_u2652_u0=and_u2643_u0&and_u2654_u0;
assign or_u740_u0=and_delayed_u65_u0|or_u739_u0;
assign and_u2653_u0=and_u2642_u0&block_GO_delayed_u42;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u65_u0<=1'h0;
else and_delayed_u65_u0<=and_u2653_u0;
end
assign and_u2654_u0=and_u2641_u0&block_GO_delayed_u42;
assign and_u2655_u0=block_GO_delayed_u42&syncEnable_u373_u0;
assign not_u553_u0=~syncEnable_u373_u0;
assign and_u2656_u0=block_GO_delayed_u42&not_u553_u0;
assign simplePinWrite_u703=and_u2657_u0&{1{and_u2657_u0}};
assign and_u2657_u0=and_u2658_u0&and_u2658_u0;
assign and_u2658_u0=and_u2659_u0&and_u2659_u0;
assign or_u741_u0=port_010c32d0_|reg_00e338d7_u0;
assign and_u2659_u0=and_u2655_u0&block_GO_delayed_u42;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00e338d7_u0<=1'h0;
else reg_00e338d7_u0<=and_u2660_u0;
end
assign and_u2660_u0=and_u2656_u0&block_GO_delayed_u42;
assign not_u554_u0=~syncEnable_u374_u0;
assign and_u2661_u0=block_GO_delayed_u42&not_u554_u0;
assign and_u2662_u0=block_GO_delayed_u42&syncEnable_u374_u0;
assign not_u555_u0=~syncEnable_u371;
assign and_u2663_u0=and_u2673_u0&syncEnable_u371;
assign and_u2664_u0=and_u2673_u0&not_u555_u0;
assign simplePinWrite_u704=and_u2665_u0&{1{and_u2665_u0}};
assign and_u2665_u0=and_u2672_u0&and_u2672_u0;
assign and_u2666_u0=and_u2670_u0&and_u2640_u0;
assign and_u2667_u0=and_u2670_u0&not_u556_u0;
assign not_u556_u0=~and_u2640_u0;
assign simplePinWrite_u705=and_u2669_u0&{1{and_u2669_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00cc41c6_u0<=1'h0;
else reg_00cc41c6_u0<=and_u2668_u0;
end
assign or_u742_u0=reg_001f57d1_u0|reg_00cc41c6_u0;
assign and_u2668_u0=and_u2667_u0&and_u2670_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_001f57d1_u0<=1'h0;
else reg_001f57d1_u0<=reg_01d1ae03_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01d1ae03_u0<=1'h0;
else reg_01d1ae03_u0<=and_u2669_u0;
end
assign and_u2669_u0=and_u2666_u0&and_u2670_u0;
assign and_u2670_u0=and_u2671_u0&and_u2671_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00f575f7_u0<=1'h0;
else reg_00f575f7_u0<=and_u2672_u0;
end
assign or_u743_u0=reg_00f575f7_u0|or_u742_u0;
assign and_u2671_u0=and_u2664_u0&and_u2673_u0;
assign and_u2672_u0=and_u2663_u0&and_u2673_u0;
assign and_u2673_u0=and_u2662_u0&block_GO_delayed_u42;
assign and_u2674_u0=and_u2661_u0&block_GO_delayed_u42;
assign or_u744_u0=or_u743_u0|and_delayed_u66_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u66_u0<=1'h0;
else and_delayed_u66_u0<=and_u2674_u0;
end
assign mux_u496=(and_u2657_u0)?1'h1:1'h0;
assign or_u745_u0=and_u2657_u0|and_u2665_u0;
assign mux_u497_u0=(and_u2645_u0)?1'h1:1'h0;
assign or_u746_u0=and_u2645_u0|and_u2657_u0;
assign doneCountIm_go_merge=simplePinWrite|simplePinWrite_u704;
assign mux_u498_u0=(and_u2645_u0)?1'h0:1'h1;
assign or_u747_u0=and_u2645_u0|and_u2665_u0;
assign scoreboard_00861902_resOr1=or_u740_u0|scoreboard_00861902_reg1;
assign scoreboard_00861902_resOr0=or_u741_u0|scoreboard_00861902_reg0;
assign bus_01994ea2_=scoreboard_00861902_and|RESET;
always @(posedge CLK)
begin
if (bus_01994ea2_)
scoreboard_00861902_reg0<=1'h0;
else if (or_u741_u0)
scoreboard_00861902_reg0<=1'h1;
else scoreboard_00861902_reg0<=scoreboard_00861902_reg0;
end
always @(posedge CLK)
begin
if (bus_01994ea2_)
scoreboard_00861902_reg2<=1'h0;
else if (or_u744_u0)
scoreboard_00861902_reg2<=1'h1;
else scoreboard_00861902_reg2<=scoreboard_00861902_reg2;
end
always @(posedge CLK)
begin
if (bus_01994ea2_)
scoreboard_00861902_reg1<=1'h0;
else if (or_u740_u0)
scoreboard_00861902_reg1<=1'h1;
else scoreboard_00861902_reg1<=scoreboard_00861902_reg1;
end
assign scoreboard_00861902_resOr2=or_u744_u0|scoreboard_00861902_reg2;
assign scoreboard_00861902_and=scoreboard_00861902_resOr0&scoreboard_00861902_resOr1&scoreboard_00861902_resOr2;
always @(posedge CLK)
begin
if (and_u2636_u0)
syncEnable_u371<=equals;
end
always @(posedge CLK)
begin
if (and_u2636_u0)
syncEnable_u372_u0<=port_0032333f_;
end
always @(posedge CLK)
begin
if (and_u2636_u0)
syncEnable_u373_u0<=port_01ce98f6_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u42<=1'h0;
else block_GO_delayed_u42<=and_u2636_u0;
end
always @(posedge CLK)
begin
if (and_u2636_u0)
syncEnable_u374_u0<=port_00c47705_;
end
always @(posedge CLK)
begin
if (and_u2636_u0)
syncEnable_u375_u0<=and_u2638_u0;
end
assign or_u748_u0=reg_0163200b_u0|scoreboard_00861902_and;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0163200b_u0<=1'h0;
else reg_0163200b_u0<=reg_0037d9b9_u0;
end
assign mux_u499_u0=(GO)?1'h0:mux_u497_u0;
assign or_u749_u0=GO|or_u746_u0;
assign mux_u500_u0=(GO)?1'h1:mux_u498_u0;
assign or_u750_u0=GO|or_u747_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0037d9b9_u0<=1'h0;
else reg_0037d9b9_u0<=GO;
end
assign or_u751_u0=GO|or_u745_u0;
assign mux_u501_u0=(GO)?1'h0:mux_u496;
assign RESULT=or_u750_u0;
assign RESULT_u1956=mux_u500_u0;
assign RESULT_u1957=or_u749_u0;
assign RESULT_u1958=mux_u499_u0;
assign RESULT_u1959=or_u751_u0;
assign RESULT_u1960=mux_u501_u0;
assign RESULT_u1961=simplePinWrite_u702;
assign RESULT_u1962=simplePinWrite_u705;
assign RESULT_u1963=simplePinWrite_u703;
assign RESULT_u1964=doneCountIm_go_merge;
assign DONE=1'h0;
endmodule



module Generation_send(CLK, RESET, GO, port_00bf371b_, port_0158b5cb_, port_00b84c6a_, port_01177a51_, port_00f76336_, port_006cd08b_, port_0197dc98_, port_0079b3b6_, RESULT, RESULT_u1965, RESULT_u1966, RESULT_u1967, RESULT_u1968, RESULT_u1969, RESULT_u1970, RESULT_u1971, RESULT_u1972, RESULT_u1973, RESULT_u1974, RESULT_u1975, RESULT_u1976, RESULT_u1977, RESULT_u1978, RESULT_u1979, RESULT_u1980, RESULT_u1981, RESULT_u1982, RESULT_u1983, RESULT_u1984, RESULT_u1985, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_00bf371b_;
input	[31:0]	port_0158b5cb_;
input		port_00b84c6a_;
input	[7:0]	port_01177a51_;
input		port_00f76336_;
input	[7:0]	port_006cd08b_;
input		port_0197dc98_;
input	[7:0]	port_0079b3b6_;
output		RESULT;
output	[31:0]	RESULT_u1965;
output		RESULT_u1966;
output	[31:0]	RESULT_u1967;
output		RESULT_u1968;
output	[31:0]	RESULT_u1969;
output	[2:0]	RESULT_u1970;
output		RESULT_u1971;
output	[31:0]	RESULT_u1972;
output	[2:0]	RESULT_u1973;
output		RESULT_u1974;
output	[31:0]	RESULT_u1975;
output	[2:0]	RESULT_u1976;
output	[15:0]	RESULT_u1977;
output	[7:0]	RESULT_u1978;
output	[7:0]	RESULT_u1979;
output		RESULT_u1980;
output	[15:0]	RESULT_u1981;
output	[7:0]	RESULT_u1982;
output	[15:0]	RESULT_u1983;
output		RESULT_u1984;
output		RESULT_u1985;
output		DONE;
wire	[31:0]	add;
wire	[31:0]	add_u1155;
wire	[31:0]	add_u1156;
wire	[31:0]	add_u1157;
wire		and_u2675_u0;
reg		done_cache_u49=1'h0;
wire		or_u752_u0;
wire	[31:0]	add_u1158;
wire	[31:0]	add_u1159;
wire	[31:0]	add_u1160;
wire	[31:0]	add_u1161;
wire		or_u753_u0;
reg		done_cache_u50_u0=1'h0;
wire		and_u2676_u0;
wire	[31:0]	add_u1162;
wire	[31:0]	add_u1163;
wire	[31:0]	add_u1164;
wire	[31:0]	add_u1165;
wire		or_u754_u0;
wire		and_u2677_u0;
reg		done_cache_u51_u0=1'h0;
wire	[31:0]	add_u1166;
wire		equals;
wire signed	[31:0]	equals_a_signed;
wire signed	[31:0]	equals_b_signed;
wire		and_u2678_u0;
wire		and_u2679_u0;
wire		not_u557_u0;
wire	[31:0]	add_u1167;
wire	[31:0]	mux_u502;
wire		and_u2680_u0;
wire		and_u2681_u0;
wire	[31:0]	mux_u503_u0;
wire	[7:0]	simplePinWrite;
wire		simplePinWrite_u706;
wire	[15:0]	simplePinWrite_u707;
wire	[7:0]	simplePinWrite_u708;
wire	[15:0]	simplePinWrite_u709;
wire		simplePinWrite_u710;
wire	[15:0]	simplePinWrite_u711;
wire	[7:0]	simplePinWrite_u712;
wire		simplePinWrite_u713;
reg	[31:0]	syncEnable_u376=32'h0;
reg		reg_00f6da00_u0=1'h0;
reg	[31:0]	syncEnable_u377_u0=32'h0;
reg		reg_00f6da00_result_delayed_u0=1'h0;
reg	[31:0]	syncEnable_u378_u0=32'h0;
assign add={port_00bf371b_[24:0], 7'b0}+{port_00bf371b_[26:0], 5'b0};
assign add_u1155={add[31:5], 5'b0}+{port_00bf371b_[27:0], 4'b0};
assign add_u1156={add_u1155[31:4], 4'b0}+port_0158b5cb_;
assign add_u1157=32'h0+add_u1156;
assign and_u2675_u0=done_cache_u49&port_0197dc98_;
always @(posedge CLK or posedge reg_00f6da00_u0 or posedge or_u752_u0)
begin
if (or_u752_u0)
done_cache_u49<=1'h0;
else if (reg_00f6da00_u0)
done_cache_u49<=1'h1;
else done_cache_u49<=done_cache_u49;
end
assign or_u752_u0=and_u2675_u0|RESET;
assign add_u1158={port_00bf371b_[24:0], 7'b0}+{port_00bf371b_[26:0], 5'b0};
assign add_u1159={add_u1158[31:5], 5'b0}+{port_00bf371b_[27:0], 4'b0};
assign add_u1160={add_u1159[31:4], 4'b0}+port_0158b5cb_;
assign add_u1161=32'h0+add_u1160;
assign or_u753_u0=and_u2676_u0|RESET;
always @(posedge CLK or posedge reg_00f6da00_u0 or posedge or_u753_u0)
begin
if (or_u753_u0)
done_cache_u50_u0<=1'h0;
else if (reg_00f6da00_u0)
done_cache_u50_u0<=1'h1;
else done_cache_u50_u0<=done_cache_u50_u0;
end
assign and_u2676_u0=done_cache_u50_u0&port_00f76336_;
assign add_u1162={port_00bf371b_[24:0], 7'b0}+{port_00bf371b_[26:0], 5'b0};
assign add_u1163={add_u1162[31:5], 5'b0}+{port_00bf371b_[27:0], 4'b0};
assign add_u1164={add_u1163[31:4], 4'b0}+port_0158b5cb_;
assign add_u1165=32'h0+add_u1164;
assign or_u754_u0=and_u2677_u0|RESET;
assign and_u2677_u0=done_cache_u51_u0&port_00b84c6a_;
always @(posedge CLK or posedge reg_00f6da00_u0 or posedge or_u754_u0)
begin
if (or_u754_u0)
done_cache_u51_u0<=1'h0;
else if (reg_00f6da00_u0)
done_cache_u51_u0<=1'h1;
else done_cache_u51_u0<=done_cache_u51_u0;
end
assign add_u1166=port_0158b5cb_+32'h1;
assign equals_a_signed=add_u1166;
assign equals_b_signed=32'hb0;
assign equals=equals_a_signed==equals_b_signed;
assign and_u2678_u0=GO&not_u557_u0;
assign and_u2679_u0=GO&equals;
assign not_u557_u0=~equals;
assign add_u1167=port_00bf371b_+32'h1;
assign mux_u502=(and_u2680_u0)?32'h0:add_u1166;
assign and_u2680_u0=and_u2679_u0&GO;
assign and_u2681_u0=and_u2678_u0&GO;
assign mux_u503_u0=(and_u2680_u0)?add_u1167:port_00bf371b_;
assign simplePinWrite=port_0079b3b6_;
assign simplePinWrite_u706=reg_00f6da00_result_delayed_u0&{1{reg_00f6da00_result_delayed_u0}};
assign simplePinWrite_u707=16'h1&{16{1'h1}};
assign simplePinWrite_u708=port_006cd08b_;
assign simplePinWrite_u709=16'h1&{16{1'h1}};
assign simplePinWrite_u710=reg_00f6da00_result_delayed_u0&{1{reg_00f6da00_result_delayed_u0}};
assign simplePinWrite_u711=16'h1&{16{1'h1}};
assign simplePinWrite_u712=port_01177a51_;
assign simplePinWrite_u713=reg_00f6da00_result_delayed_u0&{1{reg_00f6da00_result_delayed_u0}};
always @(posedge CLK)
begin
if (GO)
syncEnable_u376<=add_u1157;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00f6da00_u0<=1'h0;
else reg_00f6da00_u0<=GO;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u377_u0<=add_u1165;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00f6da00_result_delayed_u0<=1'h0;
else reg_00f6da00_result_delayed_u0<=reg_00f6da00_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u378_u0<=add_u1161;
end
assign RESULT=GO;
assign RESULT_u1965=mux_u503_u0;
assign RESULT_u1966=GO;
assign RESULT_u1967=mux_u502;
assign RESULT_u1968=reg_00f6da00_u0;
assign RESULT_u1969=syncEnable_u377_u0;
assign RESULT_u1970=3'h1;
assign RESULT_u1971=reg_00f6da00_u0;
assign RESULT_u1972=syncEnable_u378_u0;
assign RESULT_u1973=3'h1;
assign RESULT_u1974=reg_00f6da00_u0;
assign RESULT_u1975=syncEnable_u376;
assign RESULT_u1976=3'h1;
assign RESULT_u1977=simplePinWrite_u711;
assign RESULT_u1978=simplePinWrite_u708;
assign RESULT_u1979=simplePinWrite;
assign RESULT_u1980=simplePinWrite_u713;
assign RESULT_u1981=simplePinWrite_u707;
assign RESULT_u1982=simplePinWrite_u712;
assign RESULT_u1983=simplePinWrite_u709;
assign RESULT_u1984=simplePinWrite_u706;
assign RESULT_u1985=simplePinWrite_u710;
assign DONE=reg_00f6da00_result_delayed_u0;
endmodule


