// __  ___ __ ___  _ __   ___  ___ 
// \ \/ / '__/ _ \| '_ \ / _ \/ __|
//  >  <| | | (_) | | | | (_) \__ \
// /_/\_\_|  \___/|_| |_|\___/|___/
// 
// Xronos synthesizer version
// Run date: Tue 17 Nov 2015 18:39:14 +0000
// 

module Stream_to_YUV(Y_DATA, U_DATA, Y_SEND, U_ACK, V_COUNT, V_SEND, stream_ACK, U_SEND, Y_RDY, U_RDY, U_COUNT, RESET, stream_DATA, V_ACK, Y_COUNT, CLK, stream_COUNT, V_DATA, V_RDY, stream_SEND, Y_ACK);
output	[7:0]	Y_DATA;
output	[7:0]	U_DATA;
output		Y_SEND;
input		U_ACK;
wire		getPixValueU_done;
wire		getPixValueY_done;
output	[15:0]	V_COUNT;
output		V_SEND;
output		stream_ACK;
output		U_SEND;
wire		getPixValueV_go;
input		Y_RDY;
input		U_RDY;
output	[15:0]	U_COUNT;
wire		getPixValueY_go;
input		RESET;
wire		getPixValueU_go;
wire		doneCount_go;
wire		doneCount_done;
input	[7:0]	stream_DATA;
wire		getPixValueV_done;
input		V_ACK;
output	[15:0]	Y_COUNT;
input		CLK;
input	[15:0]	stream_COUNT;
output	[7:0]	V_DATA;
input		V_RDY;
input		stream_SEND;
input		Y_ACK;
wire	[7:0]	bus_019b8b17_;
wire		bus_019c80cd_;
wire		doneCount;
wire		Stream_to_YUV_doneCount_instance_DONE;
wire	[31:0]	doneCount_u12;
wire		bus_00af66a6_;
wire	[31:0]	bus_0111c215_;
wire		bus_003544db_;
wire		getPixValueU_u77;
wire	[31:0]	getPixValueU_u74;
wire		getPixValueU;
wire		Stream_to_YUV_getPixValueU_instance_DONE;
wire		getPixValueU_u73;
wire	[7:0]	getPixValueU_u75;
wire	[2:0]	getPixValueU_u76;
wire	[31:0]	getPixValueU_u72;
wire		bus_00714420_;
wire		bus_00805aeb_;
wire		bus_0109a0b9_;
wire		bus_01e4a760_;
wire	[31:0]	getPixValueY_u74;
wire	[31:0]	getPixValueY_u72;
wire		getPixValueY;
wire	[7:0]	getPixValueY_u75;
wire		Stream_to_YUV_getPixValueY_instance_DONE;
wire	[2:0]	getPixValueY_u76;
wire		getPixValueY_u73;
wire		getPixValueY_u77;
wire		bus_01538205_;
wire		scheduler_u412;
wire		scheduler_u411;
wire		scheduler_u409;
wire		scheduler_u407;
wire		scheduler_u408;
wire		scheduler_u405;
wire		scheduler;
wire		scheduler_u410;
wire		scheduler_u406;
wire		Stream_to_YUV_scheduler_instance_DONE;
wire		scheduler_u404;
wire		bus_0078d939_;
wire	[7:0]	bus_00c5d02e_;
wire	[2:0]	bus_007aaae0_;
wire		bus_010216d6_;
wire	[7:0]	bus_01af0d67_;
wire		bus_01587f61_;
wire	[31:0]	bus_004f8cb0_;
wire		bus_006b800a_;
wire	[7:0]	bus_01039998_;
wire		bus_01553d04_;
wire		getPixValueV_u126;
wire	[15:0]	getPixValueV_u128;
wire		getPixValueV_u117;
wire	[2:0]	getPixValueV_u119;
wire	[31:0]	getPixValueV_u118;
wire		getPixValueV_u131;
wire	[31:0]	getPixValueV_u116;
wire		Stream_to_YUV_getPixValueV_instance_DONE;
wire		getPixValueV_u120;
wire	[2:0]	getPixValueV_u122;
wire	[7:0]	getPixValueV_u132;
wire	[15:0]	getPixValueV_u129;
wire		getPixValueV_u123;
wire	[15:0]	getPixValueV_u127;
wire	[7:0]	getPixValueV_u125;
wire		getPixValueV;
wire	[31:0]	getPixValueV_u121;
wire	[7:0]	getPixValueV_u124;
wire		getPixValueV_u130;
wire		bus_016e3f06_;
wire		or_01a49ee9_u0;
wire		bus_00cac257_;
wire		bus_01013357_;
wire	[31:0]	bus_0015cfbb_;
wire		bus_0171e4ab_;
wire	[7:0]	bus_00d3d4db_;
wire		bus_004bebcd_;
wire		bus_00d34f5e_;
wire	[2:0]	bus_00474578_;
wire	[7:0]	bus_0053f3e6_;
assign Y_DATA=getPixValueV_u124;
assign U_DATA=getPixValueV_u125;
assign Y_SEND=getPixValueV_u130;
assign getPixValueU_done=bus_00cac257_;
assign getPixValueY_done=bus_016e3f06_;
assign V_COUNT=getPixValueV_u129;
assign V_SEND=getPixValueV_u123;
assign stream_ACK=or_01a49ee9_u0;
assign U_SEND=getPixValueV_u131;
assign getPixValueV_go=scheduler_u412;
assign U_COUNT=getPixValueV_u127;
assign getPixValueY_go=scheduler_u409;
assign getPixValueU_go=scheduler_u410;
assign doneCount_go=scheduler_u411;
assign doneCount_done=bus_00714420_;
assign getPixValueV_done=bus_00805aeb_;
assign Y_COUNT=getPixValueV_u128;
assign V_DATA=getPixValueV_u132;
Stream_to_YUV_structuralmemory_00381dd2_ Stream_to_YUV_structuralmemory_00381dd2__1(.CLK_u52(CLK), 
  .bus_00b09ec7_(bus_01e4a760_), .bus_00ae68ee_(bus_0015cfbb_), .bus_017a8cbb_(3'h1), 
  .bus_01b67484_(bus_00d34f5e_), .bus_012db760_(bus_004bebcd_), .bus_00fbddc4_(bus_00d3d4db_), 
  .bus_019b8b17_(bus_019b8b17_), .bus_019c80cd_(bus_019c80cd_));
Stream_to_YUV_doneCount Stream_to_YUV_doneCount_instance(.CLK(CLK), .RESET(bus_01e4a760_), 
  .GO(doneCount_go), .RESULT(doneCount), .RESULT_u1997(doneCount_u12), .DONE(Stream_to_YUV_doneCount_instance_DONE));
Stream_to_YUV_stateVar_state_s0 Stream_to_YUV_stateVar_state_s0_1(.bus_0149438b_(CLK), 
  .bus_00f1897f_(bus_01e4a760_), .bus_01d2957f_(scheduler), .bus_00ba0a63_(scheduler_u404), 
  .bus_00af66a6_(bus_00af66a6_));
Stream_to_YUV_stateVar_count Stream_to_YUV_stateVar_count_1(.bus_0075abd7_(CLK), 
  .bus_0164bfe0_(bus_01e4a760_), .bus_00e8137d_(getPixValueY), .bus_01f94c2f_(getPixValueY_u72), 
  .bus_013c160c_(getPixValueU), .bus_011e605c_(getPixValueU_u72), .bus_010e1bf9_(getPixValueV), 
  .bus_00d9afca_(getPixValueV_u116), .bus_01c713a7_(doneCount), .bus_001eb64b_(32'h0), 
  .bus_0111c215_(bus_0111c215_));
Stream_to_YUV_stateVar_state_s1 Stream_to_YUV_stateVar_state_s1_1(.bus_01d5eb24_(CLK), 
  .bus_0140a51f_(bus_01e4a760_), .bus_013d111b_(scheduler_u405), .bus_015b7923_(scheduler_u406), 
  .bus_003544db_(bus_003544db_));
Stream_to_YUV_getPixValueU Stream_to_YUV_getPixValueU_instance(.CLK(CLK), .RESET(bus_01e4a760_), 
  .GO(getPixValueU_go), .port_01705ac8_(bus_0111c215_), .port_00edf528_(bus_006b800a_), 
  .port_0017337e_(stream_DATA), .RESULT(getPixValueU), .RESULT_u1998(getPixValueU_u72), 
  .RESULT_u1999(getPixValueU_u73), .RESULT_u2000(getPixValueU_u74), .RESULT_u2001(getPixValueU_u75), 
  .RESULT_u2002(getPixValueU_u76), .RESULT_u2003(getPixValueU_u77), .DONE(Stream_to_YUV_getPixValueU_instance_DONE));
assign bus_00714420_=Stream_to_YUV_doneCount_instance_DONE&{1{Stream_to_YUV_doneCount_instance_DONE}};
assign bus_00805aeb_=Stream_to_YUV_getPixValueV_instance_DONE&{1{Stream_to_YUV_getPixValueV_instance_DONE}};
Stream_to_YUV_stateVar_state_s2 Stream_to_YUV_stateVar_state_s2_1(.bus_00370925_(CLK), 
  .bus_01396681_(bus_01e4a760_), .bus_0184e534_(scheduler_u407), .bus_00562eb2_(scheduler_u408), 
  .bus_0109a0b9_(bus_0109a0b9_));
Stream_to_YUV_globalreset_physical_018ec90c_ Stream_to_YUV_globalreset_physical_018ec90c__1(.bus_014bca18_(CLK), 
  .bus_01fe544c_(RESET), .bus_01e4a760_(bus_01e4a760_));
Stream_to_YUV_getPixValueY Stream_to_YUV_getPixValueY_instance(.CLK(CLK), .RESET(bus_01e4a760_), 
  .GO(getPixValueY_go), .port_01877566_(bus_0111c215_), .port_00e10874_(bus_01013357_), 
  .port_0042ccea_(stream_DATA), .RESULT(getPixValueY), .RESULT_u2004(getPixValueY_u72), 
  .RESULT_u2005(getPixValueY_u73), .RESULT_u2006(getPixValueY_u74), .RESULT_u2007(getPixValueY_u75), 
  .RESULT_u2008(getPixValueY_u76), .RESULT_u2009(getPixValueY_u77), .DONE(Stream_to_YUV_getPixValueY_instance_DONE));
Stream_to_YUV_Kicker_59 Stream_to_YUV_Kicker_59_1(.CLK(CLK), .RESET(bus_01e4a760_), 
  .bus_01538205_(bus_01538205_));
Stream_to_YUV_scheduler Stream_to_YUV_scheduler_instance(.CLK(CLK), .RESET(bus_01e4a760_), 
  .GO(bus_01538205_), .port_00ac8109_(bus_00af66a6_), .port_004cc18b_(bus_003544db_), 
  .port_01ef8e77_(bus_0109a0b9_), .port_00c1b320_(bus_0111c215_), .port_01e856ea_(getPixValueV_done), 
  .port_0002860c_(Y_RDY), .port_003a6321_(getPixValueU_done), .port_01f41769_(V_RDY), 
  .port_01e19f24_(U_RDY), .port_009dc2b3_(getPixValueY_done), .port_01060f47_(doneCount_done), 
  .port_001f0b01_(stream_SEND), .RESULT(scheduler), .RESULT_u2010(scheduler_u404), 
  .RESULT_u2011(scheduler_u405), .RESULT_u2012(scheduler_u406), .RESULT_u2013(scheduler_u407), 
  .RESULT_u2014(scheduler_u408), .RESULT_u2015(scheduler_u409), .RESULT_u2016(scheduler_u410), 
  .RESULT_u2018(scheduler_u411), .RESULT_u2017(scheduler_u412), .DONE(Stream_to_YUV_scheduler_instance_DONE));
Stream_to_YUV_simplememoryreferee_0161d552_ Stream_to_YUV_simplememoryreferee_0161d552__1(.bus_01930e79_(CLK), 
  .bus_019b487d_(bus_01e4a760_), .bus_0077fd91_(bus_01553d04_), .bus_00273fae_(bus_01039998_), 
  .bus_0035f562_(getPixValueU_u73), .bus_01208bff_(getPixValueU_u75), .bus_00599561_(getPixValueU_u74), 
  .bus_01695d49_(3'h1), .bus_01afd881_(getPixValueV_u117), .bus_00bd10ef_(getPixValueV_u118), 
  .bus_01b5288b_(3'h1), .bus_00c5d02e_(bus_00c5d02e_), .bus_004f8cb0_(bus_004f8cb0_), 
  .bus_01587f61_(bus_01587f61_), .bus_010216d6_(bus_010216d6_), .bus_007aaae0_(bus_007aaae0_), 
  .bus_006b800a_(bus_006b800a_), .bus_01af0d67_(bus_01af0d67_), .bus_0078d939_(bus_0078d939_));
Stream_to_YUV_structuralmemory_004c2570_ Stream_to_YUV_structuralmemory_004c2570__1(.CLK_u53(CLK), 
  .bus_019dd080_(bus_01e4a760_), .bus_01f84642_(bus_004f8cb0_), .bus_003b3174_(3'h1), 
  .bus_000799d1_(bus_010216d6_), .bus_01454ddc_(bus_01587f61_), .bus_00d8f36c_(bus_00c5d02e_), 
  .bus_01039998_(bus_01039998_), .bus_01553d04_(bus_01553d04_));
Stream_to_YUV_getPixValueV Stream_to_YUV_getPixValueV_instance(.CLK(CLK), .RESET(bus_01e4a760_), 
  .GO(getPixValueV_go), .port_01aef692_(bus_0111c215_), .port_01384cfe_(bus_0078d939_), 
  .port_00ab5c02_(bus_01af0d67_), .port_00af34eb_(bus_0171e4ab_), .port_004125d8_(bus_0053f3e6_), 
  .port_0097d378_(stream_DATA), .RESULT(getPixValueV), .RESULT_u2019(getPixValueV_u116), 
  .RESULT_u2020(getPixValueV_u117), .RESULT_u2021(getPixValueV_u118), .RESULT_u2022(getPixValueV_u119), 
  .RESULT_u2023(getPixValueV_u120), .RESULT_u2024(getPixValueV_u121), .RESULT_u2025(getPixValueV_u122), 
  .RESULT_u2026(getPixValueV_u123), .RESULT_u2028(getPixValueV_u124), .RESULT_u2027(getPixValueV_u125), 
  .RESULT_u2030(getPixValueV_u126), .RESULT_u2029(getPixValueV_u127), .RESULT_u2031(getPixValueV_u128), 
  .RESULT_u2032(getPixValueV_u129), .RESULT_u2033(getPixValueV_u130), .RESULT_u2035(getPixValueV_u131), 
  .RESULT_u2034(getPixValueV_u132), .DONE(Stream_to_YUV_getPixValueV_instance_DONE));
assign bus_016e3f06_=Stream_to_YUV_getPixValueY_instance_DONE&{1{Stream_to_YUV_getPixValueY_instance_DONE}};
assign or_01a49ee9_u0=getPixValueY_u77|getPixValueU_u77|getPixValueV_u126;
assign bus_00cac257_=Stream_to_YUV_getPixValueU_instance_DONE&{1{Stream_to_YUV_getPixValueU_instance_DONE}};
Stream_to_YUV_simplememoryreferee_01af975d_ Stream_to_YUV_simplememoryreferee_01af975d__1(.bus_01eef605_(CLK), 
  .bus_0159e82e_(bus_01e4a760_), .bus_01ad528e_(bus_019c80cd_), .bus_01bd925b_(bus_019b8b17_), 
  .bus_01a2b698_(getPixValueY_u73), .bus_004be9dc_(getPixValueY_u75), .bus_007ef6c2_(getPixValueY_u74), 
  .bus_004ba02e_(3'h1), .bus_00feec6d_(getPixValueV_u120), .bus_0084efad_(getPixValueV_u121), 
  .bus_00148621_(3'h1), .bus_00d3d4db_(bus_00d3d4db_), .bus_0015cfbb_(bus_0015cfbb_), 
  .bus_004bebcd_(bus_004bebcd_), .bus_00d34f5e_(bus_00d34f5e_), .bus_00474578_(bus_00474578_), 
  .bus_01013357_(bus_01013357_), .bus_0053f3e6_(bus_0053f3e6_), .bus_0171e4ab_(bus_0171e4ab_));
endmodule



module Stream_to_YUV_forge_memory_25344x8_78(CLK, EN, WE, ADDR, DIN, DOUT, DONE);
input		CLK;
input		EN;
input		WE;
input	[31:0]	ADDR;
input	[7:0]	DIN;
output	[7:0]	DOUT;
output		DONE;
wire		we_0;
wire	[7:0]	pre_dout_0;
wire		we_1;
wire	[7:0]	pre_dout_1;
reg	[7:0]	mux_out;
reg	[31:0]	ADDR_reg;
reg		wen_done;
reg		ren_done;
assign we_0=WE&(ADDR[31:14]==18'h0);
assign we_1=WE&(ADDR[31:14]==18'h1);
always @(posedge CLK)
begin
ADDR_reg<=ADDR;
end
always @(ADDR_reg or pre_dout_0 or pre_dout_1)
begin
case (ADDR_reg[31:14])18'd0:mux_out=pre_dout_0;
18'd1:mux_out=pre_dout_1;
default:mux_out=8'h0;
endcase end
always @(posedge CLK)
begin
ren_done<=EN;
wen_done<=WE;
end
assign DOUT=mux_out;
assign DONE=ren_done|wen_done;
//  Memory array element: COL: 0, ROW: 0
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_800(.CLK(CLK), .WE(we_0), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[0]), 
  .DO(pre_dout_0[0]));
//  Memory array element: COL: 0, ROW: 1
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_801(.CLK(CLK), .WE(we_0), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[1]), 
  .DO(pre_dout_0[1]));
//  Memory array element: COL: 0, ROW: 2
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_802(.CLK(CLK), .WE(we_0), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[2]), 
  .DO(pre_dout_0[2]));
//  Memory array element: COL: 0, ROW: 3
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_803(.CLK(CLK), .WE(we_0), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[3]), 
  .DO(pre_dout_0[3]));
//  Memory array element: COL: 0, ROW: 4
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_804(.CLK(CLK), .WE(we_0), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[4]), 
  .DO(pre_dout_0[4]));
//  Memory array element: COL: 0, ROW: 5
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_805(.CLK(CLK), .WE(we_0), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[5]), 
  .DO(pre_dout_0[5]));
//  Memory array element: COL: 0, ROW: 6
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_806(.CLK(CLK), .WE(we_0), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[6]), 
  .DO(pre_dout_0[6]));
//  Memory array element: COL: 0, ROW: 7
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_807(.CLK(CLK), .WE(we_0), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[7]), 
  .DO(pre_dout_0[7]));
//  Memory array element: COL: 1, ROW: 0
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_808(.CLK(CLK), .WE(we_1), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[0]), 
  .DO(pre_dout_1[0]));
//  Memory array element: COL: 1, ROW: 1
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_809(.CLK(CLK), .WE(we_1), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[1]), 
  .DO(pre_dout_1[1]));
//  Memory array element: COL: 1, ROW: 2
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_810(.CLK(CLK), .WE(we_1), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[2]), 
  .DO(pre_dout_1[2]));
//  Memory array element: COL: 1, ROW: 3
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_811(.CLK(CLK), .WE(we_1), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[3]), 
  .DO(pre_dout_1[3]));
//  Memory array element: COL: 1, ROW: 4
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_812(.CLK(CLK), .WE(we_1), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[4]), 
  .DO(pre_dout_1[4]));
//  Memory array element: COL: 1, ROW: 5
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_813(.CLK(CLK), .WE(we_1), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[5]), 
  .DO(pre_dout_1[5]));
//  Memory array element: COL: 1, ROW: 6
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_814(.CLK(CLK), .WE(we_1), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[6]), 
  .DO(pre_dout_1[6]));
//  Memory array element: COL: 1, ROW: 7
//  Initialization of Block ram now done through explicit parameter
// setting.
RAMB16_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  )RAMB16_S1_instance_815(.CLK(CLK), .WE(we_1), .EN(EN), .SSR(1'b0), .ADDR(ADDR), .DI(DIN[7]), 
  .DO(pre_dout_1[7]));
endmodule



module Stream_to_YUV_structuralmemory_00381dd2_(CLK_u52, bus_00b09ec7_, bus_00ae68ee_, bus_017a8cbb_, bus_01b67484_, bus_012db760_, bus_00fbddc4_, bus_019b8b17_, bus_019c80cd_);
input		CLK_u52;
input		bus_00b09ec7_;
input	[31:0]	bus_00ae68ee_;
input	[2:0]	bus_017a8cbb_;
input		bus_01b67484_;
input		bus_012db760_;
input	[7:0]	bus_00fbddc4_;
output	[7:0]	bus_019b8b17_;
output		bus_019c80cd_;
reg		logicalMem_1633d3c_re_delay0_u0=1'h0;
wire		or_009daac7_u0;
wire		or_008d4805_u0;
wire	[7:0]	bus_014a1fd3_;
reg		logicalMem_1633d3c_we_delay0_u0=1'h0;
always @(posedge CLK_u52 or posedge bus_00b09ec7_)
begin
if (bus_00b09ec7_)
logicalMem_1633d3c_re_delay0_u0<=1'h0;
else logicalMem_1633d3c_re_delay0_u0<=bus_01b67484_;
end
assign or_009daac7_u0=bus_01b67484_|bus_012db760_;
assign bus_019b8b17_=bus_014a1fd3_;
assign bus_019c80cd_=or_008d4805_u0;
assign or_008d4805_u0=logicalMem_1633d3c_re_delay0_u0|logicalMem_1633d3c_we_delay0_u0;
Stream_to_YUV_forge_memory_25344x8_78 Stream_to_YUV_forge_memory_25344x8_78_instance0(.CLK(CLK_u52), 
  .EN(or_009daac7_u0), .WE(bus_012db760_), .ADDR(bus_00ae68ee_), .DIN(bus_00fbddc4_), 
  .DOUT(bus_014a1fd3_), .DONE());
always @(posedge CLK_u52 or posedge bus_00b09ec7_)
begin
if (bus_00b09ec7_)
logicalMem_1633d3c_we_delay0_u0<=1'h0;
else logicalMem_1633d3c_we_delay0_u0<=bus_012db760_;
end
endmodule



module Stream_to_YUV_doneCount(CLK, RESET, GO, RESULT, RESULT_u1997, DONE);
input		CLK;
input		RESET;
input		GO;
output		RESULT;
output	[31:0]	RESULT_u1997;
output		DONE;
reg		reg_01a331ed_u0=1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01a331ed_u0<=1'h0;
else reg_01a331ed_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u1997=32'h0;
assign DONE=reg_01a331ed_u0;
endmodule



module Stream_to_YUV_stateVar_state_s0(bus_0149438b_, bus_00f1897f_, bus_01d2957f_, bus_00ba0a63_, bus_00af66a6_);
input		bus_0149438b_;
input		bus_00f1897f_;
input		bus_01d2957f_;
input		bus_00ba0a63_;
output		bus_00af66a6_;
reg		stateVar_state_s0_u35=1'h0;
assign bus_00af66a6_=stateVar_state_s0_u35;
always @(posedge bus_0149438b_ or posedge bus_00f1897f_)
begin
if (bus_00f1897f_)
stateVar_state_s0_u35<=1'h0;
else if (bus_01d2957f_)
stateVar_state_s0_u35<=bus_00ba0a63_;
end
endmodule



module Stream_to_YUV_endianswapper_006a95c8_(endianswapper_006a95c8_in, endianswapper_006a95c8_out);
input	[31:0]	endianswapper_006a95c8_in;
output	[31:0]	endianswapper_006a95c8_out;
assign endianswapper_006a95c8_out=endianswapper_006a95c8_in;
endmodule



module Stream_to_YUV_endianswapper_016b5e30_(endianswapper_016b5e30_in, endianswapper_016b5e30_out);
input	[31:0]	endianswapper_016b5e30_in;
output	[31:0]	endianswapper_016b5e30_out;
assign endianswapper_016b5e30_out=endianswapper_016b5e30_in;
endmodule



module Stream_to_YUV_stateVar_count(bus_0075abd7_, bus_0164bfe0_, bus_00e8137d_, bus_01f94c2f_, bus_013c160c_, bus_011e605c_, bus_010e1bf9_, bus_00d9afca_, bus_01c713a7_, bus_001eb64b_, bus_0111c215_);
input		bus_0075abd7_;
input		bus_0164bfe0_;
input		bus_00e8137d_;
input	[31:0]	bus_01f94c2f_;
input		bus_013c160c_;
input	[31:0]	bus_011e605c_;
input		bus_010e1bf9_;
input	[31:0]	bus_00d9afca_;
input		bus_01c713a7_;
input	[31:0]	bus_001eb64b_;
output	[31:0]	bus_0111c215_;
wire	[31:0]	endianswapper_006a95c8_out;
wire	[31:0]	endianswapper_016b5e30_out;
wire	[31:0]	mux_00bd6403_u0;
reg	[31:0]	stateVar_count_u12=32'h0;
wire		or_00fba2b0_u0;
Stream_to_YUV_endianswapper_006a95c8_ Stream_to_YUV_endianswapper_006a95c8__1(.endianswapper_006a95c8_in(stateVar_count_u12), 
  .endianswapper_006a95c8_out(endianswapper_006a95c8_out));
Stream_to_YUV_endianswapper_016b5e30_ Stream_to_YUV_endianswapper_016b5e30__1(.endianswapper_016b5e30_in(mux_00bd6403_u0), 
  .endianswapper_016b5e30_out(endianswapper_016b5e30_out));
assign mux_00bd6403_u0=({32{bus_00e8137d_}}&bus_01f94c2f_)|({32{bus_013c160c_}}&bus_011e605c_)|({32{bus_010e1bf9_}}&bus_00d9afca_)|({32{bus_01c713a7_}}&32'h0);
always @(posedge bus_0075abd7_ or posedge bus_0164bfe0_)
begin
if (bus_0164bfe0_)
stateVar_count_u12<=32'h0;
else if (or_00fba2b0_u0)
stateVar_count_u12<=endianswapper_016b5e30_out;
end
assign bus_0111c215_=endianswapper_006a95c8_out;
assign or_00fba2b0_u0=bus_00e8137d_|bus_013c160c_|bus_010e1bf9_|bus_01c713a7_;
endmodule



module Stream_to_YUV_stateVar_state_s1(bus_01d5eb24_, bus_0140a51f_, bus_013d111b_, bus_015b7923_, bus_003544db_);
input		bus_01d5eb24_;
input		bus_0140a51f_;
input		bus_013d111b_;
input		bus_015b7923_;
output		bus_003544db_;
reg		stateVar_state_s1_u35=1'h0;
assign bus_003544db_=stateVar_state_s1_u35;
always @(posedge bus_01d5eb24_ or posedge bus_0140a51f_)
begin
if (bus_0140a51f_)
stateVar_state_s1_u35<=1'h0;
else if (bus_013d111b_)
stateVar_state_s1_u35<=bus_015b7923_;
end
endmodule



module Stream_to_YUV_getPixValueU(CLK, RESET, GO, port_01705ac8_, port_00edf528_, port_0017337e_, RESULT, RESULT_u1998, RESULT_u1999, RESULT_u2000, RESULT_u2001, RESULT_u2002, RESULT_u2003, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_01705ac8_;
input		port_00edf528_;
input	[7:0]	port_0017337e_;
output		RESULT;
output	[31:0]	RESULT_u1998;
output		RESULT_u1999;
output	[31:0]	RESULT_u2000;
output	[7:0]	RESULT_u2001;
output	[2:0]	RESULT_u2002;
output		RESULT_u2003;
output		DONE;
wire		simplePinWrite;
wire	[31:0]	add;
wire		and_u2717_u0;
wire		or_u756_u0;
reg		reg_016ef135_u0=1'h0;
wire	[31:0]	add_u1190;
reg		reg_003f3515_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign add=32'h0+port_01705ac8_;
assign and_u2717_u0=reg_016ef135_u0&port_00edf528_;
assign or_u756_u0=and_u2717_u0|RESET;
always @(posedge CLK or posedge GO or posedge or_u756_u0)
begin
if (or_u756_u0)
reg_016ef135_u0<=1'h0;
else if (GO)
reg_016ef135_u0<=1'h1;
else reg_016ef135_u0<=reg_016ef135_u0;
end
assign add_u1190=port_01705ac8_+32'h1;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_003f3515_u0<=1'h0;
else reg_003f3515_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u1998=add_u1190;
assign RESULT_u1999=GO;
assign RESULT_u2000=add;
assign RESULT_u2001=port_0017337e_;
assign RESULT_u2002=3'h1;
assign RESULT_u2003=simplePinWrite;
assign DONE=reg_003f3515_u0;
endmodule



module Stream_to_YUV_stateVar_state_s2(bus_00370925_, bus_01396681_, bus_0184e534_, bus_00562eb2_, bus_0109a0b9_);
input		bus_00370925_;
input		bus_01396681_;
input		bus_0184e534_;
input		bus_00562eb2_;
output		bus_0109a0b9_;
reg		stateVar_state_s2_u33=1'h0;
always @(posedge bus_00370925_ or posedge bus_01396681_)
begin
if (bus_01396681_)
stateVar_state_s2_u33<=1'h0;
else if (bus_0184e534_)
stateVar_state_s2_u33<=bus_00562eb2_;
end
assign bus_0109a0b9_=stateVar_state_s2_u33;
endmodule



module Stream_to_YUV_globalreset_physical_018ec90c_(bus_014bca18_, bus_01fe544c_, bus_01e4a760_);
input		bus_014bca18_;
input		bus_01fe544c_;
output		bus_01e4a760_;
wire		and_01b2b09f_u0;
wire		or_00506b6d_u0;
wire		not_01abe48e_u0;
reg		final_u59=1'h1;
reg		sample_u59=1'h0;
reg		cross_u59=1'h0;
reg		glitch_u59=1'h0;
assign and_01b2b09f_u0=cross_u59&glitch_u59;
assign or_00506b6d_u0=bus_01fe544c_|final_u59;
assign not_01abe48e_u0=~and_01b2b09f_u0;
always @(posedge bus_014bca18_)
begin
final_u59<=not_01abe48e_u0;
end
always @(posedge bus_014bca18_)
begin
sample_u59<=1'h1;
end
always @(posedge bus_014bca18_)
begin
cross_u59<=sample_u59;
end
assign bus_01e4a760_=or_00506b6d_u0;
always @(posedge bus_014bca18_)
begin
glitch_u59<=cross_u59;
end
endmodule



module Stream_to_YUV_getPixValueY(CLK, RESET, GO, port_01877566_, port_00e10874_, port_0042ccea_, RESULT, RESULT_u2004, RESULT_u2005, RESULT_u2006, RESULT_u2007, RESULT_u2008, RESULT_u2009, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_01877566_;
input		port_00e10874_;
input	[7:0]	port_0042ccea_;
output		RESULT;
output	[31:0]	RESULT_u2004;
output		RESULT_u2005;
output	[31:0]	RESULT_u2006;
output	[7:0]	RESULT_u2007;
output	[2:0]	RESULT_u2008;
output		RESULT_u2009;
output		DONE;
wire		simplePinWrite;
wire	[31:0]	add;
reg		reg_016d447f_u0=1'h0;
wire		and_u2718_u0;
wire		or_u757_u0;
wire	[31:0]	add_u1191;
reg		reg_01c6f0cc_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign add=32'h0+port_01877566_;
always @(posedge CLK or posedge GO or posedge or_u757_u0)
begin
if (or_u757_u0)
reg_016d447f_u0<=1'h0;
else if (GO)
reg_016d447f_u0<=1'h1;
else reg_016d447f_u0<=reg_016d447f_u0;
end
assign and_u2718_u0=reg_016d447f_u0&port_00e10874_;
assign or_u757_u0=and_u2718_u0|RESET;
assign add_u1191=port_01877566_+32'h1;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01c6f0cc_u0<=1'h0;
else reg_01c6f0cc_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u2004=add_u1191;
assign RESULT_u2005=GO;
assign RESULT_u2006=add;
assign RESULT_u2007=port_0042ccea_;
assign RESULT_u2008=3'h1;
assign RESULT_u2009=simplePinWrite;
assign DONE=reg_01c6f0cc_u0;
endmodule



module Stream_to_YUV_Kicker_59(CLK, RESET, bus_01538205_);
input		CLK;
input		RESET;
output		bus_01538205_;
wire		bus_00359953_;
wire		bus_01b4ff55_;
wire		bus_002aae41_;
reg		kicker_res=1'h0;
wire		bus_0138d3db_;
reg		kicker_2=1'h0;
reg		kicker_1=1'h0;
assign bus_00359953_=~RESET;
assign bus_01b4ff55_=~kicker_2;
assign bus_002aae41_=bus_00359953_&kicker_1;
assign bus_01538205_=kicker_res;
always @(posedge CLK)
begin
kicker_res<=bus_0138d3db_;
end
assign bus_0138d3db_=kicker_1&bus_00359953_&bus_01b4ff55_;
always @(posedge CLK)
begin
kicker_2<=bus_002aae41_;
end
always @(posedge CLK)
begin
kicker_1<=bus_00359953_;
end
endmodule



module Stream_to_YUV_scheduler(CLK, RESET, GO, port_00ac8109_, port_004cc18b_, port_01ef8e77_, port_00c1b320_, port_01e856ea_, port_0002860c_, port_01e19f24_, port_01f41769_, port_003a6321_, port_009dc2b3_, port_01060f47_, port_001f0b01_, RESULT, RESULT_u2010, RESULT_u2011, RESULT_u2012, RESULT_u2013, RESULT_u2014, RESULT_u2015, RESULT_u2016, RESULT_u2017, RESULT_u2018, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_00ac8109_;
input		port_004cc18b_;
input		port_01ef8e77_;
input	[31:0]	port_00c1b320_;
input		port_01e856ea_;
input		port_0002860c_;
input		port_01e19f24_;
input		port_01f41769_;
input		port_003a6321_;
input		port_009dc2b3_;
input		port_01060f47_;
input		port_001f0b01_;
output		RESULT;
output		RESULT_u2010;
output		RESULT_u2011;
output		RESULT_u2012;
output		RESULT_u2013;
output		RESULT_u2014;
output		RESULT_u2015;
output		RESULT_u2016;
output		RESULT_u2017;
output		RESULT_u2018;
output		DONE;
wire		equals;
wire signed	[31:0]	equals_a_signed;
wire signed	[31:0]	equals_b_signed;
wire		and_u2719_u0;
wire		and_u2720_u0;
wire		not_u566_u0;
wire		and_u2721_u0;
wire		and_u2722_u0;
wire		and_u2723_u0;
wire		not_u567_u0;
wire		and_u2724_u0;
wire		simplePinWrite;
wire		and_u2725_u0;
wire		not_u568_u0;
wire		and_u2726_u0;
wire		and_u2727_u0;
wire		simplePinWrite_u725;
wire		and_u2728_u0;
wire		and_u2729_u0;
wire		and_u2730_u0;
wire		and_u2731_u0;
wire		and_u2732_u0;
wire		and_u2733_u0;
wire		not_u569_u0;
wire		and_u2734_u0;
wire		and_u2735_u0;
wire		and_u2736_u0;
wire		not_u570_u0;
wire		simplePinWrite_u726;
wire		and_u2737_u0;
wire		not_u571_u0;
wire		and_u2738_u0;
wire		and_u2739_u0;
wire		simplePinWrite_u727;
wire		and_u2740_u0;
wire		and_u2741_u0;
wire		and_u2742_u0;
wire		and_u2743_u0;
wire		and_u2744_u0;
wire		and_u2745_u0;
wire		not_u572_u0;
wire		and_u2746_u0;
wire		not_u573_u0;
wire		and_u2747_u0;
wire		and_u2748_u0;
wire		simplePinWrite_u728;
wire		and_u2749_u0;
wire		and_u2750_u0;
wire		and_u2751_u0;
wire		not_u574_u0;
wire		and_u2752_u0;
wire		and_u2753_u0;
wire		not_u575_u0;
wire		simplePinWrite_u729;
wire		and_u2754_u0;
wire		and_u2755_u0;
wire		and_u2756_u0;
wire		and_u2757_u0;
wire		and_u2758_u0;
wire		or_u758_u0;
wire		mux_u510;
wire		doneCount_go_merge;
wire		or_u759_u0;
wire		mux_u511_u0;
wire		mux_u512_u0;
wire		or_u760_u0;
reg		syncEnable_u379=1'h0;
reg		syncEnable_u380_u0=1'h0;
reg		syncEnable_u381_u0=1'h0;
reg		block_GO_delayed_u43=1'h0;
reg		syncEnable_u382_u0=1'h0;
reg		syncEnable_u383_u0=1'h0;
reg		syncEnable_u384_u0=1'h0;
reg		syncEnable_u385_u0=1'h0;
reg		syncEnable_u386_u0=1'h0;
reg		reg_01d006b5_u0=1'h0;
reg		reg_00b233fe_u0=1'h0;
wire		and_u2759_u0;
reg		loopControl_u43=1'h0;
reg		syncEnable_u387_u0=1'h0;
wire		or_u761_u0;
wire		mux_u513_u0;
wire		or_u762_u0;
reg		reg_01712b52_u0=1'h0;
wire		or_u763_u0;
wire		mux_u514_u0;
wire		or_u764_u0;
wire		mux_u515_u0;
reg		reg_01fd12bd_u0=1'h0;
assign equals_a_signed=port_00c1b320_;
assign equals_b_signed=32'h6300;
assign equals=equals_a_signed==equals_b_signed;
assign and_u2719_u0=port_0002860c_&port_01e19f24_;
assign and_u2720_u0=and_u2719_u0&syncEnable_u386_u0;
assign not_u566_u0=~syncEnable_u383_u0;
assign and_u2721_u0=block_GO_delayed_u43&not_u566_u0;
assign and_u2722_u0=block_GO_delayed_u43&syncEnable_u383_u0;
assign and_u2723_u0=and_u2732_u0&syncEnable_u380_u0;
assign not_u567_u0=~syncEnable_u380_u0;
assign and_u2724_u0=and_u2732_u0&not_u567_u0;
assign simplePinWrite=and_u2725_u0&{1{and_u2725_u0}};
assign and_u2725_u0=and_u2730_u0&and_u2730_u0;
assign not_u568_u0=~syncEnable_u379;
assign and_u2726_u0=and_u2731_u0&not_u568_u0;
assign and_u2727_u0=and_u2731_u0&syncEnable_u379;
assign simplePinWrite_u725=and_u2728_u0&{1{and_u2728_u0}};
assign and_u2728_u0=and_u2729_u0&and_u2729_u0;
assign and_u2729_u0=and_u2727_u0&and_u2731_u0;
assign and_u2730_u0=and_u2723_u0&and_u2732_u0;
assign and_u2731_u0=and_u2724_u0&and_u2732_u0;
assign and_u2732_u0=and_u2722_u0&block_GO_delayed_u43;
assign and_u2733_u0=block_GO_delayed_u43&not_u569_u0;
assign not_u569_u0=~syncEnable_u382_u0;
assign and_u2734_u0=block_GO_delayed_u43&syncEnable_u382_u0;
assign and_u2735_u0=and_u2744_u0&syncEnable_u380_u0;
assign and_u2736_u0=and_u2744_u0&not_u570_u0;
assign not_u570_u0=~syncEnable_u380_u0;
assign simplePinWrite_u726=and_u2737_u0&{1{and_u2737_u0}};
assign and_u2737_u0=and_u2743_u0&and_u2743_u0;
assign not_u571_u0=~syncEnable_u381_u0;
assign and_u2738_u0=and_u2742_u0&not_u571_u0;
assign and_u2739_u0=and_u2742_u0&syncEnable_u381_u0;
assign simplePinWrite_u727=and_u2740_u0&{1{and_u2740_u0}};
assign and_u2740_u0=and_u2741_u0&and_u2741_u0;
assign and_u2741_u0=and_u2739_u0&and_u2742_u0;
assign and_u2742_u0=and_u2736_u0&and_u2744_u0;
assign and_u2743_u0=and_u2735_u0&and_u2744_u0;
assign and_u2744_u0=and_u2734_u0&block_GO_delayed_u43;
assign and_u2745_u0=block_GO_delayed_u43&not_u572_u0;
assign not_u572_u0=~syncEnable_u385_u0;
assign and_u2746_u0=block_GO_delayed_u43&syncEnable_u385_u0;
assign not_u573_u0=~syncEnable_u380_u0;
assign and_u2747_u0=and_u2758_u0&not_u573_u0;
assign and_u2748_u0=and_u2758_u0&syncEnable_u380_u0;
assign simplePinWrite_u728=and_u2749_u0&{1{and_u2749_u0}};
assign and_u2749_u0=and_u2757_u0&and_u2757_u0;
assign and_u2750_u0=and_u2756_u0&not_u574_u0;
assign and_u2751_u0=and_u2756_u0&syncEnable_u384_u0;
assign not_u574_u0=~syncEnable_u384_u0;
assign and_u2752_u0=and_u2755_u0&not_u575_u0;
assign and_u2753_u0=and_u2755_u0&and_u2720_u0;
assign not_u575_u0=~and_u2720_u0;
assign simplePinWrite_u729=and_u2754_u0&{1{and_u2754_u0}};
assign and_u2754_u0=and_u2753_u0&and_u2755_u0;
assign and_u2755_u0=and_u2751_u0&and_u2756_u0;
assign and_u2756_u0=and_u2747_u0&and_u2758_u0;
assign and_u2757_u0=and_u2748_u0&and_u2758_u0;
assign and_u2758_u0=and_u2746_u0&block_GO_delayed_u43;
assign or_u758_u0=and_u2737_u0|and_u2749_u0;
assign mux_u510=(and_u2737_u0)?1'h1:1'h0;
assign doneCount_go_merge=simplePinWrite|simplePinWrite_u726|simplePinWrite_u728;
assign or_u759_u0=and_u2725_u0|and_u2737_u0;
assign mux_u511_u0=(and_u2725_u0)?1'h1:1'h0;
assign mux_u512_u0=(and_u2725_u0)?1'h0:1'h1;
assign or_u760_u0=and_u2725_u0|and_u2749_u0;
always @(posedge CLK)
begin
if (and_u2759_u0)
syncEnable_u379<=port_001f0b01_;
end
always @(posedge CLK)
begin
if (and_u2759_u0)
syncEnable_u380_u0<=equals;
end
always @(posedge CLK)
begin
if (and_u2759_u0)
syncEnable_u381_u0<=port_001f0b01_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u43<=1'h0;
else block_GO_delayed_u43<=and_u2759_u0;
end
always @(posedge CLK)
begin
if (and_u2759_u0)
syncEnable_u382_u0<=port_004cc18b_;
end
always @(posedge CLK)
begin
if (and_u2759_u0)
syncEnable_u383_u0<=port_00ac8109_;
end
always @(posedge CLK)
begin
if (and_u2759_u0)
syncEnable_u384_u0<=port_001f0b01_;
end
always @(posedge CLK)
begin
if (and_u2759_u0)
syncEnable_u385_u0<=port_01ef8e77_;
end
always @(posedge CLK)
begin
if (and_u2759_u0)
syncEnable_u386_u0<=port_01f41769_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01d006b5_u0<=1'h0;
else reg_01d006b5_u0<=reg_00b233fe_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00b233fe_u0<=1'h0;
else reg_00b233fe_u0<=and_u2759_u0;
end
assign and_u2759_u0=or_u761_u0&or_u761_u0;
always @(posedge CLK or posedge syncEnable_u387_u0)
begin
if (syncEnable_u387_u0)
loopControl_u43<=1'h0;
else loopControl_u43<=reg_01d006b5_u0;
end
always @(posedge CLK)
begin
if (reg_01712b52_u0)
syncEnable_u387_u0<=RESET;
end
assign or_u761_u0=loopControl_u43|reg_01712b52_u0;
assign mux_u513_u0=(GO)?1'h0:mux_u511_u0;
assign or_u762_u0=GO|or_u759_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01712b52_u0<=1'h0;
else reg_01712b52_u0<=reg_01fd12bd_u0;
end
assign or_u763_u0=GO|or_u760_u0;
assign mux_u514_u0=(GO)?1'h1:mux_u512_u0;
assign or_u764_u0=GO|or_u758_u0;
assign mux_u515_u0=(GO)?1'h0:mux_u510;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01fd12bd_u0<=1'h0;
else reg_01fd12bd_u0<=GO;
end
assign RESULT=or_u763_u0;
assign RESULT_u2010=mux_u514_u0;
assign RESULT_u2011=or_u762_u0;
assign RESULT_u2012=mux_u513_u0;
assign RESULT_u2013=or_u764_u0;
assign RESULT_u2014=mux_u515_u0;
assign RESULT_u2015=simplePinWrite_u725;
assign RESULT_u2016=simplePinWrite_u727;
assign RESULT_u2017=simplePinWrite_u729;
assign RESULT_u2018=doneCount_go_merge;
assign DONE=1'h0;
endmodule



module Stream_to_YUV_simplememoryreferee_0161d552_(bus_01930e79_, bus_019b487d_, bus_0077fd91_, bus_00273fae_, bus_0035f562_, bus_01208bff_, bus_00599561_, bus_01695d49_, bus_01afd881_, bus_00bd10ef_, bus_01b5288b_, bus_00c5d02e_, bus_004f8cb0_, bus_01587f61_, bus_010216d6_, bus_007aaae0_, bus_006b800a_, bus_01af0d67_, bus_0078d939_);
input		bus_01930e79_;
input		bus_019b487d_;
input		bus_0077fd91_;
input	[7:0]	bus_00273fae_;
input		bus_0035f562_;
input	[7:0]	bus_01208bff_;
input	[31:0]	bus_00599561_;
input	[2:0]	bus_01695d49_;
input		bus_01afd881_;
input	[31:0]	bus_00bd10ef_;
input	[2:0]	bus_01b5288b_;
output	[7:0]	bus_00c5d02e_;
output	[31:0]	bus_004f8cb0_;
output		bus_01587f61_;
output		bus_010216d6_;
output	[2:0]	bus_007aaae0_;
output		bus_006b800a_;
output	[7:0]	bus_01af0d67_;
output		bus_0078d939_;
wire	[31:0]	mux_00fc8151_u0;
wire	[7:0]	mux_01beb1c2_u0;
wire		and_00f8e2a3_u0;
wire		or_00e4f7c0_u0;
wire		not_014d4d8d_u0;
reg		done_qual_u156=1'h0;
wire		not_01dc431a_u0;
wire		and_01fea0ef_u0;
wire		or_00828814_u0;
wire		or_01c8a78d_u0;
reg		done_qual_u157_u0=1'h0;
assign mux_00fc8151_u0=(bus_0035f562_)?bus_00599561_:bus_00bd10ef_;
assign mux_01beb1c2_u0=({8{bus_0035f562_}}&bus_01208bff_);
assign and_00f8e2a3_u0=or_00828814_u0&bus_0077fd91_;
assign or_00e4f7c0_u0=bus_0035f562_|done_qual_u157_u0;
assign not_014d4d8d_u0=~bus_0077fd91_;
always @(posedge bus_01930e79_)
begin
if (bus_019b487d_)
done_qual_u156<=1'h0;
else done_qual_u156<=bus_01afd881_;
end
assign not_01dc431a_u0=~bus_0077fd91_;
assign and_01fea0ef_u0=or_00e4f7c0_u0&bus_0077fd91_;
assign or_00828814_u0=bus_01afd881_|done_qual_u156;
assign bus_00c5d02e_=mux_01beb1c2_u0;
assign bus_004f8cb0_=mux_00fc8151_u0;
assign bus_01587f61_=bus_0035f562_;
assign bus_010216d6_=or_01c8a78d_u0;
assign bus_007aaae0_=3'h1;
assign bus_006b800a_=and_01fea0ef_u0;
assign bus_01af0d67_=bus_00273fae_;
assign bus_0078d939_=and_00f8e2a3_u0;
assign or_01c8a78d_u0=bus_0035f562_|bus_01afd881_;
always @(posedge bus_01930e79_)
begin
if (bus_019b487d_)
done_qual_u157_u0<=1'h0;
else done_qual_u157_u0<=bus_0035f562_;
end
endmodule



module Stream_to_YUV_structuralmemory_004c2570_(CLK_u53, bus_019dd080_, bus_01f84642_, bus_003b3174_, bus_000799d1_, bus_01454ddc_, bus_00d8f36c_, bus_01039998_, bus_01553d04_);
input		CLK_u53;
input		bus_019dd080_;
input	[31:0]	bus_01f84642_;
input	[2:0]	bus_003b3174_;
input		bus_000799d1_;
input		bus_01454ddc_;
input	[7:0]	bus_00d8f36c_;
output	[7:0]	bus_01039998_;
output		bus_01553d04_;
reg		logicalMem_d8f2a6_we_delay0_u0=1'h0;
reg		logicalMem_d8f2a6_re_delay0_u0=1'h0;
wire		or_0055b9f9_u0;
wire		or_01c57902_u0;
wire	[7:0]	bus_00d16f44_;
always @(posedge CLK_u53 or posedge bus_019dd080_)
begin
if (bus_019dd080_)
logicalMem_d8f2a6_we_delay0_u0<=1'h0;
else logicalMem_d8f2a6_we_delay0_u0<=bus_01454ddc_;
end
always @(posedge CLK_u53 or posedge bus_019dd080_)
begin
if (bus_019dd080_)
logicalMem_d8f2a6_re_delay0_u0<=1'h0;
else logicalMem_d8f2a6_re_delay0_u0<=bus_000799d1_;
end
assign or_0055b9f9_u0=bus_000799d1_|bus_01454ddc_;
assign bus_01039998_=bus_00d16f44_;
assign bus_01553d04_=or_01c57902_u0;
assign or_01c57902_u0=logicalMem_d8f2a6_re_delay0_u0|logicalMem_d8f2a6_we_delay0_u0;
Stream_to_YUV_forge_memory_25344x8_78 Stream_to_YUV_forge_memory_25344x8_78_instance1(.CLK(CLK_u53), 
  .EN(or_0055b9f9_u0), .WE(bus_01454ddc_), .ADDR(bus_01f84642_), .DIN(bus_00d8f36c_), 
  .DOUT(bus_00d16f44_), .DONE());
endmodule



module Stream_to_YUV_getPixValueV(CLK, RESET, GO, port_01aef692_, port_01384cfe_, port_00ab5c02_, port_00af34eb_, port_004125d8_, port_0097d378_, RESULT, RESULT_u2019, RESULT_u2020, RESULT_u2021, RESULT_u2022, RESULT_u2023, RESULT_u2024, RESULT_u2025, RESULT_u2026, RESULT_u2027, RESULT_u2028, RESULT_u2029, RESULT_u2030, RESULT_u2031, RESULT_u2032, RESULT_u2033, RESULT_u2034, RESULT_u2035, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_01aef692_;
input		port_01384cfe_;
input	[7:0]	port_00ab5c02_;
input		port_00af34eb_;
input	[7:0]	port_004125d8_;
input	[7:0]	port_0097d378_;
output		RESULT;
output	[31:0]	RESULT_u2019;
output		RESULT_u2020;
output	[31:0]	RESULT_u2021;
output	[2:0]	RESULT_u2022;
output		RESULT_u2023;
output	[31:0]	RESULT_u2024;
output	[2:0]	RESULT_u2025;
output		RESULT_u2026;
output	[7:0]	RESULT_u2027;
output	[7:0]	RESULT_u2028;
output	[15:0]	RESULT_u2029;
output		RESULT_u2030;
output	[15:0]	RESULT_u2031;
output	[15:0]	RESULT_u2032;
output		RESULT_u2033;
output	[7:0]	RESULT_u2034;
output		RESULT_u2035;
output		DONE;
wire		simplePinWrite;
wire	[31:0]	add;
reg		done_cache_u52=1'h0;
wire		or_u765_u0;
wire		and_u2760_u0;
wire	[31:0]	add_u1192;
reg		done_cache_u53_u0=1'h0;
wire		or_u766_u0;
wire		and_u2761_u0;
wire	[31:0]	add_u1193;
wire		simplePinWrite_u730;
wire	[7:0]	simplePinWrite_u731;
wire	[15:0]	simplePinWrite_u732;
wire		simplePinWrite_u733;
wire	[7:0]	simplePinWrite_u734;
wire	[15:0]	simplePinWrite_u735;
wire		simplePinWrite_u736;
wire	[7:0]	simplePinWrite_u737;
wire	[15:0]	simplePinWrite_u738;
reg		reg_0109c23b_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign add=32'h0+port_01aef692_;
always @(posedge CLK or posedge GO or posedge or_u765_u0)
begin
if (or_u765_u0)
done_cache_u52<=1'h0;
else if (GO)
done_cache_u52<=1'h1;
else done_cache_u52<=done_cache_u52;
end
assign or_u765_u0=and_u2760_u0|RESET;
assign and_u2760_u0=done_cache_u52&port_00af34eb_;
assign add_u1192=32'h0+port_01aef692_;
always @(posedge CLK or posedge GO or posedge or_u766_u0)
begin
if (or_u766_u0)
done_cache_u53_u0<=1'h0;
else if (GO)
done_cache_u53_u0<=1'h1;
else done_cache_u53_u0<=done_cache_u53_u0;
end
assign or_u766_u0=and_u2761_u0|RESET;
assign and_u2761_u0=done_cache_u53_u0&port_01384cfe_;
assign add_u1193=port_01aef692_+32'h1;
assign simplePinWrite_u730=reg_0109c23b_u0&{1{reg_0109c23b_u0}};
assign simplePinWrite_u731=port_004125d8_;
assign simplePinWrite_u732=16'h1&{16{1'h1}};
assign simplePinWrite_u733=reg_0109c23b_u0&{1{reg_0109c23b_u0}};
assign simplePinWrite_u734=port_00ab5c02_;
assign simplePinWrite_u735=16'h1&{16{1'h1}};
assign simplePinWrite_u736=GO&{1{GO}};
assign simplePinWrite_u737=port_0097d378_;
assign simplePinWrite_u738=16'h1&{16{1'h1}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0109c23b_u0<=1'h0;
else reg_0109c23b_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u2019=add_u1193;
assign RESULT_u2020=GO;
assign RESULT_u2021=add_u1192;
assign RESULT_u2022=3'h1;
assign RESULT_u2023=GO;
assign RESULT_u2024=add;
assign RESULT_u2025=3'h1;
assign RESULT_u2026=simplePinWrite_u736;
assign RESULT_u2027=simplePinWrite_u734;
assign RESULT_u2028=simplePinWrite_u731;
assign RESULT_u2029=simplePinWrite_u735;
assign RESULT_u2030=simplePinWrite;
assign RESULT_u2031=simplePinWrite_u732;
assign RESULT_u2032=simplePinWrite_u738;
assign RESULT_u2033=simplePinWrite_u730;
assign RESULT_u2034=simplePinWrite_u737;
assign RESULT_u2035=simplePinWrite_u733;
assign DONE=reg_0109c23b_u0;
endmodule



module Stream_to_YUV_simplememoryreferee_01af975d_(bus_01eef605_, bus_0159e82e_, bus_01ad528e_, bus_01bd925b_, bus_01a2b698_, bus_004be9dc_, bus_007ef6c2_, bus_004ba02e_, bus_00feec6d_, bus_0084efad_, bus_00148621_, bus_00d3d4db_, bus_0015cfbb_, bus_004bebcd_, bus_00d34f5e_, bus_00474578_, bus_01013357_, bus_0053f3e6_, bus_0171e4ab_);
input		bus_01eef605_;
input		bus_0159e82e_;
input		bus_01ad528e_;
input	[7:0]	bus_01bd925b_;
input		bus_01a2b698_;
input	[7:0]	bus_004be9dc_;
input	[31:0]	bus_007ef6c2_;
input	[2:0]	bus_004ba02e_;
input		bus_00feec6d_;
input	[31:0]	bus_0084efad_;
input	[2:0]	bus_00148621_;
output	[7:0]	bus_00d3d4db_;
output	[31:0]	bus_0015cfbb_;
output		bus_004bebcd_;
output		bus_00d34f5e_;
output	[2:0]	bus_00474578_;
output		bus_01013357_;
output	[7:0]	bus_0053f3e6_;
output		bus_0171e4ab_;
wire		not_0176e40a_u0;
wire	[31:0]	mux_00b839bf_u0;
wire		and_00bb81d2_u0;
reg		done_qual_u158_u0=1'h0;
wire	[7:0]	mux_0135dad2_u0;
wire		or_018bd378_u0;
wire		and_01fa47f8_u0;
wire		not_00ca1355_u0;
reg		done_qual_u159_u0=1'h0;
wire		or_010f4a8a_u0;
wire		or_015c5808_u0;
assign bus_00d3d4db_=mux_0135dad2_u0;
assign bus_0015cfbb_=mux_00b839bf_u0;
assign bus_004bebcd_=bus_01a2b698_;
assign bus_00d34f5e_=or_015c5808_u0;
assign bus_00474578_=3'h1;
assign bus_01013357_=and_01fa47f8_u0;
assign bus_0053f3e6_=bus_01bd925b_;
assign bus_0171e4ab_=and_00bb81d2_u0;
assign not_0176e40a_u0=~bus_01ad528e_;
assign mux_00b839bf_u0=(bus_01a2b698_)?bus_007ef6c2_:bus_0084efad_;
assign and_00bb81d2_u0=or_010f4a8a_u0&bus_01ad528e_;
always @(posedge bus_01eef605_)
begin
if (bus_0159e82e_)
done_qual_u158_u0<=1'h0;
else done_qual_u158_u0<=bus_01a2b698_;
end
assign mux_0135dad2_u0=({8{bus_01a2b698_}}&bus_004be9dc_);
assign or_018bd378_u0=bus_01a2b698_|done_qual_u158_u0;
assign and_01fa47f8_u0=or_018bd378_u0&bus_01ad528e_;
assign not_00ca1355_u0=~bus_01ad528e_;
always @(posedge bus_01eef605_)
begin
if (bus_0159e82e_)
done_qual_u159_u0<=1'h0;
else done_qual_u159_u0<=bus_00feec6d_;
end
assign or_010f4a8a_u0=bus_00feec6d_|done_qual_u159_u0;
assign or_015c5808_u0=bus_01a2b698_|bus_00feec6d_;
endmodule


