// __  ___ __ ___  _ __   ___  ___ 
// \ \/ / '__/ _ \| '_ \ / _ \/ __|
//  >  <| | | (_) | | | | (_) \__ \
// /_/\_\_|  \___/|_| |_|\___/|___/
// 
// Xronos synthesizer version
// Run date: Tue 17 Nov 2015 16:03:58 +0000
// 

module PROCESS(Bout_DATA, RESET, Gout_SEND, Gout_DATA, Gin_DATA, Gin_COUNT, Rout_DATA, Rin_SEND, Bin_DATA, Gin_ACK, Rout_ACK, Bin_ACK, Gin_SEND, Bin_SEND, Bout_ACK, Rin_COUNT, CLK, Rout_COUNT, Gout_COUNT, Bin_COUNT, Bout_RDY, Rout_SEND, Gout_ACK, Rin_ACK, Bout_COUNT, Rin_DATA, Bout_SEND, Gout_RDY, Rout_RDY);
wire		doneCountIm_done;
output	[7:0]	Bout_DATA;
input		RESET;
wire		doneCountIm_go;
output		Gout_SEND;
output	[7:0]	Gout_DATA;
input	[7:0]	Gin_DATA;
input	[15:0]	Gin_COUNT;
output	[7:0]	Rout_DATA;
input		Rin_SEND;
input	[7:0]	Bin_DATA;
wire		send_go;
output		Gin_ACK;
wire		drawRectangle_done;
input		Rout_ACK;
output		Bin_ACK;
wire		getValueRGB_go;
input		Gin_SEND;
input		Bin_SEND;
input		Bout_ACK;
wire		send_done;
input	[15:0]	Rin_COUNT;
wire		getValueRGB_done;
input		CLK;
output	[15:0]	Rout_COUNT;
output	[15:0]	Gout_COUNT;
input	[15:0]	Bin_COUNT;
input		Bout_RDY;
output		Rout_SEND;
input		Gout_ACK;
wire		drawRectangle_go;
output		Rin_ACK;
output	[15:0]	Bout_COUNT;
input	[7:0]	Rin_DATA;
output		Bout_SEND;
input		Gout_RDY;
input		Rout_RDY;
wire		bus_01cbaafe_;
wire		bus_01a55e8c_;
wire	[7:0]	bus_01253f88_;
wire	[31:0]	doneCountIm_u4;
wire		PROCESS_doneCountIm_instance_DONE;
wire		doneCountIm;
wire		bus_01f7d5fe_;
wire		bus_00e248e8_;
wire	[7:0]	bus_01abaecf_;
wire		bus_00c4ebf0_;
wire		bus_00a49847_;
wire	[31:0]	bus_00b4b9d0_;
wire		bus_01047a38_;
wire		bus_00f0c433_;
wire	[7:0]	bus_00e37882_;
wire	[2:0]	bus_00e765a2_;
wire		bus_0153aeef_;
wire		bus_01292474_;
wire		bus_00e6429a_;
wire	[7:0]	bus_01e84f7c_;
wire		bus_019dab71_;
wire	[2:0]	bus_01754a4a_;
wire		bus_0194c9bb_;
wire	[31:0]	bus_01dfb2dc_;
wire		bus_01493d37_;
wire	[7:0]	bus_018c4737_;
wire	[31:0]	bus_0011e612_;
wire		bus_018e3bd5_;
wire		bus_01ff0a92_;
wire	[31:0]	bus_0120c5dc_;
wire		bus_00d6ed62_;
wire	[7:0]	bus_01a38a4e_;
wire		bus_000fcc00_;
wire		bus_00c9542f_;
wire	[7:0]	bus_01140234_;
wire	[2:0]	bus_00414afd_;
wire		scheduler_u234;
wire		scheduler_u235;
wire		scheduler_u233;
wire		scheduler;
wire		scheduler_u237;
wire		scheduler_u232;
wire		scheduler_u240;
wire		scheduler_u238;
wire		PROCESS_scheduler_instance_DONE;
wire		scheduler_u236;
wire		scheduler_u239;
wire		bus_008e2aa8_;
wire	[7:0]	bus_019151a3_;
wire		bus_010aabe7_;
wire		bus_010cc662_;
wire	[31:0]	drawRectangle_u100;
wire	[7:0]	drawRectangle_u93;
wire	[31:0]	drawRectangle_u112;
wire		drawRectangle_u99;
wire		drawRectangle;
wire		PROCESS_drawRectangle_instance_DONE;
wire	[2:0]	drawRectangle_u106;
wire	[2:0]	drawRectangle_u110;
wire		drawRectangle_u95;
wire	[31:0]	drawRectangle_u104;
wire	[7:0]	drawRectangle_u113;
wire	[31:0]	drawRectangle_u108;
wire	[2:0]	drawRectangle_u114;
wire	[7:0]	drawRectangle_u105;
wire	[31:0]	drawRectangle_u96;
wire		drawRectangle_u111;
wire	[2:0]	drawRectangle_u98;
wire		drawRectangle_u107;
wire	[2:0]	drawRectangle_u102;
wire	[7:0]	drawRectangle_u97;
wire	[7:0]	drawRectangle_u109;
wire	[7:0]	drawRectangle_u101;
wire	[2:0]	drawRectangle_u94;
wire		drawRectangle_u103;
wire	[31:0]	drawRectangle_u92;
wire	[15:0]	send_u132;
wire	[7:0]	send_u131;
wire	[2:0]	send_u120;
wire		send_u129;
wire		send_u121;
wire	[2:0]	send_u117;
wire	[31:0]	send_u122;
wire	[2:0]	send_u123;
wire		send_u118;
wire		send_u130;
wire	[7:0]	send_u127;
wire		PROCESS_send_instance_DONE;
wire	[15:0]	send_u125;
wire	[15:0]	send_u126;
wire		send_u128;
wire	[31:0]	send_u112;
wire	[31:0]	send_u119;
wire	[31:0]	send_u116;
wire		send_u113;
wire	[7:0]	send_u124;
wire		send;
wire	[31:0]	send_u114;
wire		send_u115;
wire		bus_0001e8b0_;
wire		bus_01726b76_;
wire		PROCESS_getValueRGB_instance_DONE;
wire		getValueRGB_u88;
wire	[31:0]	getValueRGB_u72;
wire		getValueRGB_u89;
wire	[2:0]	getValueRGB_u78;
wire	[2:0]	getValueRGB_u82;
wire		getValueRGB;
wire	[7:0]	getValueRGB_u77;
wire		getValueRGB_u83;
wire	[31:0]	getValueRGB_u84;
wire		getValueRGB_u73;
wire		getValueRGB_u79;
wire	[2:0]	getValueRGB_u86;
wire		getValueRGB_u75;
wire		getValueRGB_u87;
wire	[7:0]	getValueRGB_u85;
wire	[31:0]	getValueRGB_u76;
wire	[31:0]	getValueRGB_u74;
wire	[31:0]	getValueRGB_u80;
wire	[7:0]	getValueRGB_u81;
wire		bus_010a585d_;
wire		bus_014f17a8_;
wire	[31:0]	bus_01a2f21a_;
wire	[7:0]	bus_00f11bd2_;
wire		bus_01a2e3de_;
wire	[2:0]	bus_017fc3a3_;
wire		bus_00a7282d_;
wire		bus_00e30286_;
wire	[2:0]	bus_015b67b7_;
wire	[31:0]	bus_013b413c_;
wire		bus_0166f79c_;
wire	[7:0]	bus_01154382_;
wire		bus_00709018_;
wire		bus_013a80a2_;
wire		bus_01a77aad_;
wire		bus_0088e767_;
wire	[31:0]	bus_009f3313_;
wire		bus_0174247e_;
wire		bus_0160b5ac_;
wire		bus_01ba61a9_;
wire	[2:0]	bus_001f0d05_;
wire	[7:0]	bus_005e8c9d_;
wire	[31:0]	bus_00a07c46_;
wire		bus_00ebe0d9_;
wire	[7:0]	bus_009a9712_;
wire		bus_010bfe43_;
assign doneCountIm_done=bus_008e2aa8_;
assign Bout_DATA=send_u127;
assign doneCountIm_go=scheduler_u238;
assign Gout_SEND=send_u129;
assign Gout_DATA=send_u131;
assign Rout_DATA=send_u124;
assign send_go=scheduler_u237;
assign Gin_ACK=getValueRGB_u87;
assign drawRectangle_done=bus_0153aeef_;
assign Bin_ACK=getValueRGB_u88;
assign getValueRGB_go=scheduler_u240;
assign send_done=bus_01f7d5fe_;
assign getValueRGB_done=bus_01a77aad_;
assign Rout_COUNT=send_u125;
assign Gout_COUNT=send_u126;
assign Rout_SEND=send_u128;
assign drawRectangle_go=scheduler_u239;
assign Rin_ACK=getValueRGB_u89;
assign Bout_COUNT=send_u132;
assign Bout_SEND=send_u130;
PROCESS_structuralmemory_007e03a9_ PROCESS_structuralmemory_007e03a9__1(.CLK_u16(CLK), 
  .bus_01e9149a_(bus_01726b76_), .bus_012d2ddd_(bus_00b4b9d0_), .bus_00d10fdb_(3'h1), 
  .bus_00368442_(bus_01047a38_), .bus_0085b9f1_(bus_00e248e8_), .bus_00052497_(bus_00e37882_), 
  .bus_01265ced_(bus_00a07c46_), .bus_0161b4b5_(3'h1), .bus_01ee8bcf_(bus_01ba61a9_), 
  .bus_01cc8379_(8'h0), .bus_01253f88_(bus_01253f88_), .bus_01a55e8c_(bus_01a55e8c_), 
  .bus_01cbaafe_(bus_01cbaafe_));
PROCESS_doneCountIm PROCESS_doneCountIm_instance(.CLK(CLK), .RESET(bus_01726b76_), 
  .GO(doneCountIm_go), .RESULT(doneCountIm), .RESULT_u974(doneCountIm_u4), .DONE(PROCESS_doneCountIm_instance_DONE));
assign bus_01f7d5fe_=PROCESS_send_instance_DONE&{1{PROCESS_send_instance_DONE}};
PROCESS_simplememoryreferee_0168d4ac_ PROCESS_simplememoryreferee_0168d4ac__1(.bus_002efc6b_(CLK), 
  .bus_00bdf4b1_(bus_01726b76_), .bus_00726ac2_(bus_01a55e8c_), .bus_01d05e5e_(bus_01253f88_), 
  .bus_0129fa02_(getValueRGB_u83), .bus_0116c937_(getValueRGB_u85), .bus_01e4689a_(getValueRGB_u84), 
  .bus_017f1f8e_(3'h1), .bus_00db3f63_(drawRectangle_u107), .bus_016ac854_(8'h0), 
  .bus_015e547b_(drawRectangle_u108), .bus_000c420f_(3'h1), .bus_00524eae_(send_u118), 
  .bus_00b948fb_(send_u119), .bus_00b85ff8_(3'h1), .bus_00e37882_(bus_00e37882_), 
  .bus_00b4b9d0_(bus_00b4b9d0_), .bus_00e248e8_(bus_00e248e8_), .bus_01047a38_(bus_01047a38_), 
  .bus_00e765a2_(bus_00e765a2_), .bus_00f0c433_(bus_00f0c433_), .bus_00c4ebf0_(bus_00c4ebf0_), 
  .bus_01abaecf_(bus_01abaecf_), .bus_00a49847_(bus_00a49847_));
assign bus_0153aeef_=PROCESS_drawRectangle_instance_DONE&{1{PROCESS_drawRectangle_instance_DONE}};
PROCESS_simplememoryreferee_008d75ed_ PROCESS_simplememoryreferee_008d75ed__1(.bus_008d58e2_(CLK), 
  .bus_01c667f8_(bus_01726b76_), .bus_00cbc4cb_(bus_010cc662_), .bus_0000b302_(bus_019151a3_), 
  .bus_006ddb3e_(getValueRGB_u75), .bus_0114ac01_(getValueRGB_u77), .bus_00abe46b_(getValueRGB_u76), 
  .bus_0192fda0_(3'h1), .bus_018b18c7_(drawRectangle_u111), .bus_006ceacc_(8'h0), 
  .bus_0042fe7f_(drawRectangle_u112), .bus_01ebf7fd_(3'h1), .bus_010dbf54_(send_u115), 
  .bus_01493a7a_(send_u116), .bus_00c1b626_(3'h1), .bus_01e84f7c_(bus_01e84f7c_), 
  .bus_01dfb2dc_(bus_01dfb2dc_), .bus_01292474_(bus_01292474_), .bus_0194c9bb_(bus_0194c9bb_), 
  .bus_01754a4a_(bus_01754a4a_), .bus_01493d37_(bus_01493d37_), .bus_00e6429a_(bus_00e6429a_), 
  .bus_018c4737_(bus_018c4737_), .bus_019dab71_(bus_019dab71_));
PROCESS_stateVar_count_x PROCESS_stateVar_count_x_1(.bus_019f1881_(CLK), .bus_0001ca4b_(bus_01726b76_), 
  .bus_01e587c8_(getValueRGB), .bus_01a62129_(getValueRGB_u72), .bus_018dcccc_(doneCountIm), 
  .bus_01fdaab8_(32'h0), .bus_00ec91dd_(send), .bus_00e1da25_(send_u112), .bus_0011e612_(bus_0011e612_));
PROCESS_simplememoryreferee_00574fd0_ PROCESS_simplememoryreferee_00574fd0__1(.bus_00a2ffed_(CLK), 
  .bus_01506088_(bus_01726b76_), .bus_0046cd71_(bus_00ebe0d9_), .bus_01e7134a_(bus_009a9712_), 
  .bus_01ab54eb_(getValueRGB_u79), .bus_019de908_(getValueRGB_u81), .bus_00eeb7ef_(getValueRGB_u80), 
  .bus_01bb6b7e_(3'h1), .bus_0144f414_(drawRectangle), .bus_01fd78d5_(8'hff), .bus_00fee334_(drawRectangle_u92), 
  .bus_019a14f9_(3'h1), .bus_01a25756_(send_u121), .bus_003ad8b6_(send_u122), .bus_01085033_(3'h1), 
  .bus_01a38a4e_(bus_01a38a4e_), .bus_0120c5dc_(bus_0120c5dc_), .bus_01ff0a92_(bus_01ff0a92_), 
  .bus_000fcc00_(bus_000fcc00_), .bus_00414afd_(bus_00414afd_), .bus_018e3bd5_(bus_018e3bd5_), 
  .bus_00d6ed62_(bus_00d6ed62_), .bus_01140234_(bus_01140234_), .bus_00c9542f_(bus_00c9542f_));
PROCESS_scheduler PROCESS_scheduler_instance(.CLK(CLK), .RESET(bus_01726b76_), 
  .GO(bus_00709018_), .port_0182596d_(bus_013a80a2_), .port_0148d67c_(bus_0001e8b0_), 
  .port_015a802e_(bus_0088e767_), .port_01ead277_(bus_0011e612_), .port_0041cb2b_(Bout_RDY), 
  .port_00082475_(Bin_SEND), .port_00795ad5_(Rin_SEND), .port_01ac2e8e_(doneCountIm_done), 
  .port_0059f665_(send_done), .port_01c6ea35_(getValueRGB_done), .port_008097c7_(Gout_RDY), 
  .port_017d6741_(Rout_RDY), .port_0195d97b_(drawRectangle_done), .port_012cd222_(Gin_SEND), 
  .RESULT(scheduler), .RESULT_u975(scheduler_u232), .RESULT_u976(scheduler_u233), 
  .RESULT_u977(scheduler_u234), .RESULT_u978(scheduler_u235), .RESULT_u979(scheduler_u236), 
  .RESULT_u980(scheduler_u237), .RESULT_u982(scheduler_u238), .RESULT_u981(scheduler_u239), 
  .RESULT_u983(scheduler_u240), .DONE(PROCESS_scheduler_instance_DONE));
assign bus_008e2aa8_=PROCESS_doneCountIm_instance_DONE&{1{PROCESS_doneCountIm_instance_DONE}};
PROCESS_structuralmemory_00814577_ PROCESS_structuralmemory_00814577__1(.CLK_u17(CLK), 
  .bus_01c52148_(bus_01726b76_), .bus_00890cb8_(bus_01dfb2dc_), .bus_014efb86_(3'h1), 
  .bus_00aef9ca_(bus_0194c9bb_), .bus_00e5479e_(bus_01292474_), .bus_010d9e31_(bus_01e84f7c_), 
  .bus_0000f23b_(bus_013b413c_), .bus_00b89a1d_(3'h1), .bus_01d3fa4a_(bus_0166f79c_), 
  .bus_0118cc44_(8'h0), .bus_019151a3_(bus_019151a3_), .bus_010cc662_(bus_010cc662_), 
  .bus_010aabe7_(bus_010aabe7_));
PROCESS_drawRectangle PROCESS_drawRectangle_instance(.CLK(CLK), .RESET(bus_01726b76_), 
  .GO(drawRectangle_go), .port_006015e8_(bus_00d6ed62_), .port_01cb501c_(bus_014f17a8_), 
  .port_00e850d8_(bus_0160b5ac_), .port_014d58fd_(bus_00a7282d_), .port_0130bfa1_(bus_00c4ebf0_), 
  .port_01243a78_(bus_00e6429a_), .RESULT_u991(drawRectangle), .RESULT_u992(drawRectangle_u92), 
  .RESULT_u993(drawRectangle_u93), .RESULT_u994(drawRectangle_u94), .RESULT_u999(drawRectangle_u95), 
  .RESULT_u1000(drawRectangle_u96), .RESULT_u1001(drawRectangle_u97), .RESULT_u1002(drawRectangle_u98), 
  .RESULT_u1003(drawRectangle_u99), .RESULT_u1004(drawRectangle_u100), .RESULT_u1005(drawRectangle_u101), 
  .RESULT_u1006(drawRectangle_u102), .RESULT_u995(drawRectangle_u103), .RESULT_u996(drawRectangle_u104), 
  .RESULT_u997(drawRectangle_u105), .RESULT_u998(drawRectangle_u106), .RESULT(drawRectangle_u107), 
  .RESULT_u984(drawRectangle_u108), .RESULT_u985(drawRectangle_u109), .RESULT_u986(drawRectangle_u110), 
  .RESULT_u987(drawRectangle_u111), .RESULT_u988(drawRectangle_u112), .RESULT_u989(drawRectangle_u113), 
  .RESULT_u990(drawRectangle_u114), .DONE(PROCESS_drawRectangle_instance_DONE));
PROCESS_send PROCESS_send_instance(.CLK(CLK), .RESET(bus_01726b76_), .GO(send_go), 
  .port_01245fcb_(bus_0011e612_), .port_00c7b822_(bus_009f3313_), .port_010e3311_(bus_019dab71_), 
  .port_0148441b_(bus_018c4737_), .port_00817c5e_(bus_00a49847_), .port_015914f6_(bus_01abaecf_), 
  .port_012755fe_(bus_00c9542f_), .port_0041b215_(bus_01140234_), .RESULT(send), 
  .RESULT_u1007(send_u112), .RESULT_u1008(send_u113), .RESULT_u1009(send_u114), 
  .RESULT_u1013(send_u115), .RESULT_u1014(send_u116), .RESULT_u1015(send_u117), 
  .RESULT_u1010(send_u118), .RESULT_u1011(send_u119), .RESULT_u1012(send_u120), 
  .RESULT_u1016(send_u121), .RESULT_u1017(send_u122), .RESULT_u1018(send_u123), 
  .RESULT_u1019(send_u124), .RESULT_u1020(send_u125), .RESULT_u1021(send_u126), 
  .RESULT_u1022(send_u127), .RESULT_u1023(send_u128), .RESULT_u1025(send_u129), 
  .RESULT_u1024(send_u130), .RESULT_u1027(send_u131), .RESULT_u1026(send_u132), 
  .DONE(PROCESS_send_instance_DONE));
PROCESS_stateVar_state_s1 PROCESS_stateVar_state_s1_1(.bus_0008ca2f_(CLK), .bus_0111fdbc_(bus_01726b76_), 
  .bus_00e044d2_(scheduler_u233), .bus_01b1cd40_(scheduler_u234), .bus_0001e8b0_(bus_0001e8b0_));
PROCESS_globalreset_physical_016c3655_ PROCESS_globalreset_physical_016c3655__1(.bus_00046cea_(CLK), 
  .bus_010f4e6e_(RESET), .bus_01726b76_(bus_01726b76_));
PROCESS_getValueRGB PROCESS_getValueRGB_instance(.CLK(CLK), .RESET(bus_01726b76_), 
  .GO(getValueRGB_go), .port_00285e4f_(bus_0011e612_), .port_00028fcf_(bus_009f3313_), 
  .port_00100350_(bus_01493d37_), .port_01f41dbb_(bus_018e3bd5_), .port_00612b21_(bus_00f0c433_), 
  .port_0011132f_(Bin_DATA), .port_00b6c0b7_(Rin_DATA), .port_003f6d63_(Gin_DATA), 
  .RESULT(getValueRGB), .RESULT_u1028(getValueRGB_u72), .RESULT_u1029(getValueRGB_u73), 
  .RESULT_u1030(getValueRGB_u74), .RESULT_u1035(getValueRGB_u75), .RESULT_u1036(getValueRGB_u76), 
  .RESULT_u1037(getValueRGB_u77), .RESULT_u1038(getValueRGB_u78), .RESULT_u1039(getValueRGB_u79), 
  .RESULT_u1040(getValueRGB_u80), .RESULT_u1041(getValueRGB_u81), .RESULT_u1042(getValueRGB_u82), 
  .RESULT_u1031(getValueRGB_u83), .RESULT_u1032(getValueRGB_u84), .RESULT_u1033(getValueRGB_u85), 
  .RESULT_u1034(getValueRGB_u86), .RESULT_u1043(getValueRGB_u87), .RESULT_u1044(getValueRGB_u88), 
  .RESULT_u1045(getValueRGB_u89), .DONE(PROCESS_getValueRGB_instance_DONE));
PROCESS_simplememoryreferee_018cecb6_ PROCESS_simplememoryreferee_018cecb6__1(.bus_004bdde8_(CLK), 
  .bus_00d5e4f7_(bus_01726b76_), .bus_0074cb0b_(bus_010bfe43_), .bus_0092b9ff_(8'h0), 
  .bus_01655295_(drawRectangle_u95), .bus_00ba52c3_(8'hff), .bus_0092895d_(drawRectangle_u96), 
  .bus_0018d135_(3'h1), .bus_00f11bd2_(bus_00f11bd2_), .bus_01a2f21a_(bus_01a2f21a_), 
  .bus_010a585d_(bus_010a585d_), .bus_01a2e3de_(bus_01a2e3de_), .bus_017fc3a3_(bus_017fc3a3_), 
  .bus_014f17a8_(bus_014f17a8_));
PROCESS_simplememoryreferee_01df3566_ PROCESS_simplememoryreferee_01df3566__1(.bus_00f883fe_(CLK), 
  .bus_01a1d096_(bus_01726b76_), .bus_01662e30_(bus_010aabe7_), .bus_018b8df6_(8'h0), 
  .bus_006e6d0c_(drawRectangle_u103), .bus_00cc16ec_(8'h0), .bus_00dda92a_(drawRectangle_u104), 
  .bus_00381fab_(3'h1), .bus_01154382_(bus_01154382_), .bus_013b413c_(bus_013b413c_), 
  .bus_0166f79c_(bus_0166f79c_), .bus_00e30286_(bus_00e30286_), .bus_015b67b7_(bus_015b67b7_), 
  .bus_00a7282d_(bus_00a7282d_));
PROCESS_Kicker_34 PROCESS_Kicker_34_1(.CLK(CLK), .RESET(bus_01726b76_), .bus_00709018_(bus_00709018_));
PROCESS_stateVar_state_s0 PROCESS_stateVar_state_s0_1(.bus_01ae46ae_(CLK), .bus_00a25ac8_(bus_01726b76_), 
  .bus_000bdb25_(scheduler), .bus_0045f0e9_(scheduler_u232), .bus_013a80a2_(bus_013a80a2_));
assign bus_01a77aad_=PROCESS_getValueRGB_instance_DONE&{1{PROCESS_getValueRGB_instance_DONE}};
PROCESS_stateVar_state_s2 PROCESS_stateVar_state_s2_1(.bus_01855671_(CLK), .bus_00ee2f23_(bus_01726b76_), 
  .bus_01cf20d2_(scheduler_u235), .bus_01948536_(scheduler_u236), .bus_0088e767_(bus_0088e767_));
PROCESS_stateVar_count_y PROCESS_stateVar_count_y_1(.bus_01722449_(CLK), .bus_00ac4f02_(bus_01726b76_), 
  .bus_01303bc0_(getValueRGB_u73), .bus_01483acc_(getValueRGB_u74), .bus_0047b12a_(send_u113), 
  .bus_01c6542c_(send_u114), .bus_009f3313_(bus_009f3313_));
PROCESS_simplememoryreferee_01e963df_ PROCESS_simplememoryreferee_01e963df__1(.bus_00eb96d7_(CLK), 
  .bus_00fc372b_(bus_01726b76_), .bus_0123c590_(bus_01cbaafe_), .bus_00395682_(8'h0), 
  .bus_007262df_(drawRectangle_u99), .bus_00577cfe_(8'h0), .bus_004fde95_(drawRectangle_u100), 
  .bus_01289d14_(3'h1), .bus_005e8c9d_(bus_005e8c9d_), .bus_00a07c46_(bus_00a07c46_), 
  .bus_01ba61a9_(bus_01ba61a9_), .bus_0174247e_(bus_0174247e_), .bus_001f0d05_(bus_001f0d05_), 
  .bus_0160b5ac_(bus_0160b5ac_));
PROCESS_structuralmemory_0145fced_ PROCESS_structuralmemory_0145fced__1(.CLK_u18(CLK), 
  .bus_00ecf8c6_(bus_01726b76_), .bus_00703654_(bus_0120c5dc_), .bus_002a587c_(3'h1), 
  .bus_012a3f30_(bus_000fcc00_), .bus_00a4b4e9_(bus_01ff0a92_), .bus_01e65d20_(bus_01a38a4e_), 
  .bus_00dfcb52_(bus_01a2f21a_), .bus_00d32323_(3'h1), .bus_00681dd1_(bus_010a585d_), 
  .bus_006d22dd_(8'hff), .bus_009a9712_(bus_009a9712_), .bus_00ebe0d9_(bus_00ebe0d9_), 
  .bus_010bfe43_(bus_010bfe43_));
endmodule



module PROCESS_forge_memory_25344x8_27(CLK, ENA, WEA, DINA, ENB, WEB, DINB, ADDRA, ADDRB, DOUTA, DONEA, DONEB);
input		CLK;
input		ENA;
input		WEA;
input	[7:0]	DINA;
input		ENB;
input		WEB;
input	[7:0]	DINB;
input	[31:0]	ADDRA;
input	[31:0]	ADDRB;
output	[7:0]	DOUTA;
output		DONEA;
output		DONEB;
wire		wea_0;
wire		web_0;
wire	[7:0]	pre_douta_0;
wire		wea_1;
wire		web_1;
wire	[7:0]	pre_douta_1;
reg	[7:0]	mux_outa;
reg	[31:0]	ADDRA_reg;
reg	[31:0]	ADDRB_reg;
reg	[7:0]	mux_outb;
wire	[7:0]	pre_doutb_0;
wire	[7:0]	pre_doutb_1;
reg		rea_done;
reg		web_done;
reg		wea_done;
assign wea_0=WEA&(ADDRA[31:14]==18'h0);
assign web_0=WEB&(ADDRB[31:14]==18'h0);
assign wea_1=WEA&(ADDRA[31:14]==18'h1);
assign web_1=WEB&(ADDRB[31:14]==18'h1);
always @(posedge CLK)
begin
ADDRA_reg<=ADDRA;
end
always @(ADDRA_reg or pre_douta_0 or pre_douta_1)
begin
case (ADDRA_reg[31:14])18'd0:mux_outa=pre_douta_0;
18'd1:mux_outa=pre_douta_1;
default:mux_outa=8'h0;
endcase end
always @(posedge CLK)
begin
ADDRB_reg<=ADDRB;
end
always @(ADDRB_reg or pre_doutb_0 or pre_doutb_1)
begin
case (ADDRB_reg[31:14])18'd0:mux_outb=pre_doutb_0;
18'd1:mux_outb=pre_doutb_1;
default:mux_outb=8'h0;
endcase end
always @(posedge CLK)
begin
wea_done<=WEA;
rea_done<=ENA;
web_done<=WEB;
end
assign DONEA=wea_done|rea_done;
assign DONEB=web_done;
assign DOUTA=mux_outa;
// Memory array element: COL: 0, ROW: 0
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_64(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[0]), .DOA(pre_douta_0[0]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[0]), .DOB());
// Memory array element: COL: 0, ROW: 1
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_65(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[1]), .DOA(pre_douta_0[1]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[1]), .DOB());
// Memory array element: COL: 0, ROW: 2
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_66(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[2]), .DOA(pre_douta_0[2]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[2]), .DOB());
// Memory array element: COL: 0, ROW: 3
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_67(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[3]), .DOA(pre_douta_0[3]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[3]), .DOB());
// Memory array element: COL: 0, ROW: 4
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_68(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[4]), .DOA(pre_douta_0[4]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[4]), .DOB());
// Memory array element: COL: 0, ROW: 5
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_69(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[5]), .DOA(pre_douta_0[5]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[5]), .DOB());
// Memory array element: COL: 0, ROW: 6
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_70(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[6]), .DOA(pre_douta_0[6]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[6]), .DOB());
// Memory array element: COL: 0, ROW: 7
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_71(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[7]), .DOA(pre_douta_0[7]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[7]), .DOB());
// Memory array element: COL: 1, ROW: 0
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_72(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[0]), .DOA(pre_douta_1[0]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[0]), .DOB());
// Memory array element: COL: 1, ROW: 1
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_73(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[1]), .DOA(pre_douta_1[1]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[1]), .DOB());
// Memory array element: COL: 1, ROW: 2
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_74(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[2]), .DOA(pre_douta_1[2]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[2]), .DOB());
// Memory array element: COL: 1, ROW: 3
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_75(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[3]), .DOA(pre_douta_1[3]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[3]), .DOB());
// Memory array element: COL: 1, ROW: 4
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_76(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[4]), .DOA(pre_douta_1[4]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[4]), .DOB());
// Memory array element: COL: 1, ROW: 5
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_77(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[5]), .DOA(pre_douta_1[5]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[5]), .DOB());
// Memory array element: COL: 1, ROW: 6
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_78(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[6]), .DOA(pre_douta_1[6]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[6]), .DOB());
// Memory array element: COL: 1, ROW: 7
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_79(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[7]), .DOA(pre_douta_1[7]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[7]), .DOB());
endmodule



module PROCESS_structuralmemory_007e03a9_(CLK_u16, bus_01e9149a_, bus_012d2ddd_, bus_00d10fdb_, bus_00368442_, bus_0085b9f1_, bus_00052497_, bus_01265ced_, bus_0161b4b5_, bus_01ee8bcf_, bus_01cc8379_, bus_01253f88_, bus_01a55e8c_, bus_01cbaafe_);
input		CLK_u16;
input		bus_01e9149a_;
input	[31:0]	bus_012d2ddd_;
input	[2:0]	bus_00d10fdb_;
input		bus_00368442_;
input		bus_0085b9f1_;
input	[7:0]	bus_00052497_;
input	[31:0]	bus_01265ced_;
input	[2:0]	bus_0161b4b5_;
input		bus_01ee8bcf_;
input	[7:0]	bus_01cc8379_;
output	[7:0]	bus_01253f88_;
output		bus_01a55e8c_;
output		bus_01cbaafe_;
wire		or_00c21277_u0;
reg		logicalMem_532106_we_delay0_u0=1'h0;
wire		or_009b6252_u0;
wire	[7:0]	bus_0175a1a1_;
reg		logicalMem_532106_re_delay0_u0=1'h0;
reg		logicalMem_532106_we_delay0_u1_u0=1'h0;
assign or_00c21277_u0=bus_00368442_|bus_0085b9f1_;
always @(posedge CLK_u16 or posedge bus_01e9149a_)
begin
if (bus_01e9149a_)
logicalMem_532106_we_delay0_u0<=1'h0;
else logicalMem_532106_we_delay0_u0<=bus_01ee8bcf_;
end
assign or_009b6252_u0=logicalMem_532106_re_delay0_u0|logicalMem_532106_we_delay0_u1_u0;
PROCESS_forge_memory_25344x8_27 PROCESS_forge_memory_25344x8_27_instance0(.CLK(CLK_u16), 
  .ENA(or_00c21277_u0), .WEA(bus_0085b9f1_), .DINA(bus_00052497_), .ADDRA(bus_012d2ddd_), 
  .DOUTA(bus_0175a1a1_), .DONEA(), .ENB(bus_01ee8bcf_), .WEB(bus_01ee8bcf_), .DINB(8'h0), 
  .ADDRB(bus_01265ced_), .DONEB());
always @(posedge CLK_u16 or posedge bus_01e9149a_)
begin
if (bus_01e9149a_)
logicalMem_532106_re_delay0_u0<=1'h0;
else logicalMem_532106_re_delay0_u0<=bus_00368442_;
end
always @(posedge CLK_u16 or posedge bus_01e9149a_)
begin
if (bus_01e9149a_)
logicalMem_532106_we_delay0_u1_u0<=1'h0;
else logicalMem_532106_we_delay0_u1_u0<=bus_0085b9f1_;
end
assign bus_01253f88_=bus_0175a1a1_;
assign bus_01a55e8c_=or_009b6252_u0;
assign bus_01cbaafe_=logicalMem_532106_we_delay0_u0;
endmodule



module PROCESS_doneCountIm(CLK, RESET, GO, RESULT, RESULT_u974, DONE);
input		CLK;
input		RESET;
input		GO;
output		RESULT;
output	[31:0]	RESULT_u974;
output		DONE;
reg		reg_01b28dd2_u0=1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01b28dd2_u0<=1'h0;
else reg_01b28dd2_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u974=32'h0;
assign DONE=reg_01b28dd2_u0;
endmodule



module PROCESS_simplememoryreferee_0168d4ac_(bus_002efc6b_, bus_00bdf4b1_, bus_00726ac2_, bus_01d05e5e_, bus_0129fa02_, bus_0116c937_, bus_01e4689a_, bus_017f1f8e_, bus_00db3f63_, bus_016ac854_, bus_015e547b_, bus_000c420f_, bus_00524eae_, bus_00b948fb_, bus_00b85ff8_, bus_00e37882_, bus_00b4b9d0_, bus_00e248e8_, bus_01047a38_, bus_00e765a2_, bus_00f0c433_, bus_00c4ebf0_, bus_01abaecf_, bus_00a49847_);
input		bus_002efc6b_;
input		bus_00bdf4b1_;
input		bus_00726ac2_;
input	[7:0]	bus_01d05e5e_;
input		bus_0129fa02_;
input	[7:0]	bus_0116c937_;
input	[31:0]	bus_01e4689a_;
input	[2:0]	bus_017f1f8e_;
input		bus_00db3f63_;
input	[7:0]	bus_016ac854_;
input	[31:0]	bus_015e547b_;
input	[2:0]	bus_000c420f_;
input		bus_00524eae_;
input	[31:0]	bus_00b948fb_;
input	[2:0]	bus_00b85ff8_;
output	[7:0]	bus_00e37882_;
output	[31:0]	bus_00b4b9d0_;
output		bus_00e248e8_;
output		bus_01047a38_;
output	[2:0]	bus_00e765a2_;
output		bus_00f0c433_;
output		bus_00c4ebf0_;
output	[7:0]	bus_01abaecf_;
output		bus_00a49847_;
wire		or_01dcc1eb_u0;
reg		done_qual_u52=1'h0;
wire		not_0116e714_u0;
reg		done_qual_u53_u0=1'h0;
wire		not_00e2a673_u0;
wire		or_000cfd82_u0;
wire		and_00178c33_u0;
wire		or_008a84d9_u0;
wire		not_006b23c2_u0;
wire		and_012c9613_u0;
wire		or_007be30b_u0;
wire		or_00e5647d_u0;
wire	[31:0]	mux_01b88a32_u0;
reg		done_qual_u54_u0=1'h0;
wire	[7:0]	mux_0125a345_u0;
wire		and_01a9e64e_u0;
assign or_01dcc1eb_u0=bus_0129fa02_|bus_00db3f63_;
always @(posedge bus_002efc6b_)
begin
if (bus_00bdf4b1_)
done_qual_u52<=1'h0;
else done_qual_u52<=bus_0129fa02_;
end
assign not_0116e714_u0=~bus_00726ac2_;
always @(posedge bus_002efc6b_)
begin
if (bus_00bdf4b1_)
done_qual_u53_u0<=1'h0;
else done_qual_u53_u0<=bus_00524eae_;
end
assign not_00e2a673_u0=~bus_00726ac2_;
assign or_000cfd82_u0=bus_00db3f63_|done_qual_u54_u0;
assign and_00178c33_u0=or_000cfd82_u0&bus_00726ac2_;
assign bus_00e37882_=mux_0125a345_u0;
assign bus_00b4b9d0_=mux_01b88a32_u0;
assign bus_00e248e8_=or_01dcc1eb_u0;
assign bus_01047a38_=or_007be30b_u0;
assign bus_00e765a2_=3'h1;
assign bus_00f0c433_=and_01a9e64e_u0;
assign bus_00c4ebf0_=and_00178c33_u0;
assign bus_01abaecf_=bus_01d05e5e_;
assign bus_00a49847_=and_012c9613_u0;
assign or_008a84d9_u0=bus_00524eae_|done_qual_u53_u0;
assign not_006b23c2_u0=~bus_00726ac2_;
assign and_012c9613_u0=or_008a84d9_u0&bus_00726ac2_;
assign or_007be30b_u0=bus_0129fa02_|bus_00db3f63_|bus_00524eae_;
assign or_00e5647d_u0=bus_0129fa02_|done_qual_u52;
assign mux_01b88a32_u0=({32{bus_0129fa02_}}&bus_01e4689a_)|({32{bus_00db3f63_}}&bus_015e547b_)|({32{bus_00524eae_}}&bus_00b948fb_);
always @(posedge bus_002efc6b_)
begin
if (bus_00bdf4b1_)
done_qual_u54_u0<=1'h0;
else done_qual_u54_u0<=bus_00db3f63_;
end
assign mux_0125a345_u0=(bus_0129fa02_)?bus_0116c937_:8'h0;
assign and_01a9e64e_u0=or_00e5647d_u0&bus_00726ac2_;
endmodule



module PROCESS_simplememoryreferee_008d75ed_(bus_008d58e2_, bus_01c667f8_, bus_00cbc4cb_, bus_0000b302_, bus_006ddb3e_, bus_0114ac01_, bus_00abe46b_, bus_0192fda0_, bus_018b18c7_, bus_006ceacc_, bus_0042fe7f_, bus_01ebf7fd_, bus_010dbf54_, bus_01493a7a_, bus_00c1b626_, bus_01e84f7c_, bus_01dfb2dc_, bus_01292474_, bus_0194c9bb_, bus_01754a4a_, bus_01493d37_, bus_00e6429a_, bus_018c4737_, bus_019dab71_);
input		bus_008d58e2_;
input		bus_01c667f8_;
input		bus_00cbc4cb_;
input	[7:0]	bus_0000b302_;
input		bus_006ddb3e_;
input	[7:0]	bus_0114ac01_;
input	[31:0]	bus_00abe46b_;
input	[2:0]	bus_0192fda0_;
input		bus_018b18c7_;
input	[7:0]	bus_006ceacc_;
input	[31:0]	bus_0042fe7f_;
input	[2:0]	bus_01ebf7fd_;
input		bus_010dbf54_;
input	[31:0]	bus_01493a7a_;
input	[2:0]	bus_00c1b626_;
output	[7:0]	bus_01e84f7c_;
output	[31:0]	bus_01dfb2dc_;
output		bus_01292474_;
output		bus_0194c9bb_;
output	[2:0]	bus_01754a4a_;
output		bus_01493d37_;
output		bus_00e6429a_;
output	[7:0]	bus_018c4737_;
output		bus_019dab71_;
wire	[7:0]	mux_005ded21_u0;
wire		and_00992a01_u0;
reg		done_qual_u55_u0=1'h0;
wire		or_01475a54_u0;
wire		or_010e156c_u0;
wire		and_00ce4cdb_u0;
wire		or_00cb99d8_u0;
wire		and_00d9087a_u0;
wire		not_01830537_u0;
wire		or_001970f7_u0;
wire		not_0122a79f_u0;
wire	[31:0]	mux_01598a57_u0;
wire		not_0074a570_u0;
reg		done_qual_u56_u0=1'h0;
reg		done_qual_u57_u0=1'h0;
wire		or_0031b077_u0;
assign mux_005ded21_u0=(bus_006ddb3e_)?bus_0114ac01_:8'h0;
assign and_00992a01_u0=or_00cb99d8_u0&bus_00cbc4cb_;
always @(posedge bus_008d58e2_)
begin
if (bus_01c667f8_)
done_qual_u55_u0<=1'h0;
else done_qual_u55_u0<=bus_010dbf54_;
end
assign bus_01e84f7c_=mux_005ded21_u0;
assign bus_01dfb2dc_=mux_01598a57_u0;
assign bus_01292474_=or_01475a54_u0;
assign bus_0194c9bb_=or_010e156c_u0;
assign bus_01754a4a_=3'h1;
assign bus_01493d37_=and_00992a01_u0;
assign bus_00e6429a_=and_00d9087a_u0;
assign bus_018c4737_=bus_0000b302_;
assign bus_019dab71_=and_00ce4cdb_u0;
assign or_01475a54_u0=bus_006ddb3e_|bus_018b18c7_;
assign or_010e156c_u0=bus_006ddb3e_|bus_018b18c7_|bus_010dbf54_;
assign and_00ce4cdb_u0=or_001970f7_u0&bus_00cbc4cb_;
assign or_00cb99d8_u0=bus_006ddb3e_|done_qual_u56_u0;
assign and_00d9087a_u0=or_0031b077_u0&bus_00cbc4cb_;
assign not_01830537_u0=~bus_00cbc4cb_;
assign or_001970f7_u0=bus_010dbf54_|done_qual_u55_u0;
assign not_0122a79f_u0=~bus_00cbc4cb_;
assign mux_01598a57_u0=({32{bus_006ddb3e_}}&bus_00abe46b_)|({32{bus_018b18c7_}}&bus_0042fe7f_)|({32{bus_010dbf54_}}&bus_01493a7a_);
assign not_0074a570_u0=~bus_00cbc4cb_;
always @(posedge bus_008d58e2_)
begin
if (bus_01c667f8_)
done_qual_u56_u0<=1'h0;
else done_qual_u56_u0<=bus_006ddb3e_;
end
always @(posedge bus_008d58e2_)
begin
if (bus_01c667f8_)
done_qual_u57_u0<=1'h0;
else done_qual_u57_u0<=bus_018b18c7_;
end
assign or_0031b077_u0=bus_018b18c7_|done_qual_u57_u0;
endmodule



module PROCESS_endianswapper_00494325_(endianswapper_00494325_in, endianswapper_00494325_out);
input	[31:0]	endianswapper_00494325_in;
output	[31:0]	endianswapper_00494325_out;
assign endianswapper_00494325_out=endianswapper_00494325_in;
endmodule



module PROCESS_endianswapper_00a457a0_(endianswapper_00a457a0_in, endianswapper_00a457a0_out);
input	[31:0]	endianswapper_00a457a0_in;
output	[31:0]	endianswapper_00a457a0_out;
assign endianswapper_00a457a0_out=endianswapper_00a457a0_in;
endmodule



module PROCESS_stateVar_count_x(bus_019f1881_, bus_0001ca4b_, bus_01e587c8_, bus_01a62129_, bus_018dcccc_, bus_01fdaab8_, bus_00ec91dd_, bus_00e1da25_, bus_0011e612_);
input		bus_019f1881_;
input		bus_0001ca4b_;
input		bus_01e587c8_;
input	[31:0]	bus_01a62129_;
input		bus_018dcccc_;
input	[31:0]	bus_01fdaab8_;
input		bus_00ec91dd_;
input	[31:0]	bus_00e1da25_;
output	[31:0]	bus_0011e612_;
wire	[31:0]	endianswapper_00494325_out;
wire		or_00d283d5_u0;
wire	[31:0]	mux_008d0206_u0;
wire	[31:0]	endianswapper_00a457a0_out;
reg	[31:0]	stateVar_count_x_u4=32'h0;
PROCESS_endianswapper_00494325_ PROCESS_endianswapper_00494325__1(.endianswapper_00494325_in(mux_008d0206_u0), 
  .endianswapper_00494325_out(endianswapper_00494325_out));
assign or_00d283d5_u0=bus_01e587c8_|bus_018dcccc_|bus_00ec91dd_;
assign mux_008d0206_u0=({32{bus_01e587c8_}}&bus_01a62129_)|({32{bus_018dcccc_}}&32'h0)|({32{bus_00ec91dd_}}&bus_00e1da25_);
assign bus_0011e612_=endianswapper_00a457a0_out;
PROCESS_endianswapper_00a457a0_ PROCESS_endianswapper_00a457a0__1(.endianswapper_00a457a0_in(stateVar_count_x_u4), 
  .endianswapper_00a457a0_out(endianswapper_00a457a0_out));
always @(posedge bus_019f1881_ or posedge bus_0001ca4b_)
begin
if (bus_0001ca4b_)
stateVar_count_x_u4<=32'h0;
else if (or_00d283d5_u0)
stateVar_count_x_u4<=endianswapper_00494325_out;
end
endmodule



module PROCESS_simplememoryreferee_00574fd0_(bus_00a2ffed_, bus_01506088_, bus_0046cd71_, bus_01e7134a_, bus_01ab54eb_, bus_019de908_, bus_00eeb7ef_, bus_01bb6b7e_, bus_0144f414_, bus_01fd78d5_, bus_00fee334_, bus_019a14f9_, bus_01a25756_, bus_003ad8b6_, bus_01085033_, bus_01a38a4e_, bus_0120c5dc_, bus_01ff0a92_, bus_000fcc00_, bus_00414afd_, bus_018e3bd5_, bus_00d6ed62_, bus_01140234_, bus_00c9542f_);
input		bus_00a2ffed_;
input		bus_01506088_;
input		bus_0046cd71_;
input	[7:0]	bus_01e7134a_;
input		bus_01ab54eb_;
input	[7:0]	bus_019de908_;
input	[31:0]	bus_00eeb7ef_;
input	[2:0]	bus_01bb6b7e_;
input		bus_0144f414_;
input	[7:0]	bus_01fd78d5_;
input	[31:0]	bus_00fee334_;
input	[2:0]	bus_019a14f9_;
input		bus_01a25756_;
input	[31:0]	bus_003ad8b6_;
input	[2:0]	bus_01085033_;
output	[7:0]	bus_01a38a4e_;
output	[31:0]	bus_0120c5dc_;
output		bus_01ff0a92_;
output		bus_000fcc00_;
output	[2:0]	bus_00414afd_;
output		bus_018e3bd5_;
output		bus_00d6ed62_;
output	[7:0]	bus_01140234_;
output		bus_00c9542f_;
wire		or_016121b0_u0;
wire		or_011934bb_u0;
reg		done_qual_u58_u0=1'h0;
reg		done_qual_u59_u0=1'h0;
wire		and_012777dd_u0;
wire		and_00b20115_u0;
wire		not_01137431_u0;
wire		and_0190910c_u0;
reg		done_qual_u60_u0=1'h0;
wire	[7:0]	mux_01d6032b_u0;
wire		or_00278af0_u0;
wire		or_019749b6_u0;
wire		not_003da544_u0;
wire	[31:0]	mux_00427167_u0;
wire		not_0149a6f6_u0;
wire		or_008914da_u0;
assign or_016121b0_u0=bus_01a25756_|done_qual_u58_u0;
assign or_011934bb_u0=bus_0144f414_|done_qual_u59_u0;
always @(posedge bus_00a2ffed_)
begin
if (bus_01506088_)
done_qual_u58_u0<=1'h0;
else done_qual_u58_u0<=bus_01a25756_;
end
always @(posedge bus_00a2ffed_)
begin
if (bus_01506088_)
done_qual_u59_u0<=1'h0;
else done_qual_u59_u0<=bus_0144f414_;
end
assign and_012777dd_u0=or_00278af0_u0&bus_0046cd71_;
assign and_00b20115_u0=or_016121b0_u0&bus_0046cd71_;
assign not_01137431_u0=~bus_0046cd71_;
assign and_0190910c_u0=or_011934bb_u0&bus_0046cd71_;
always @(posedge bus_00a2ffed_)
begin
if (bus_01506088_)
done_qual_u60_u0<=1'h0;
else done_qual_u60_u0<=bus_01ab54eb_;
end
assign mux_01d6032b_u0=(bus_01ab54eb_)?bus_019de908_:8'hff;
assign bus_01a38a4e_=mux_01d6032b_u0;
assign bus_0120c5dc_=mux_00427167_u0;
assign bus_01ff0a92_=or_008914da_u0;
assign bus_000fcc00_=or_019749b6_u0;
assign bus_00414afd_=3'h1;
assign bus_018e3bd5_=and_012777dd_u0;
assign bus_00d6ed62_=and_0190910c_u0;
assign bus_01140234_=bus_01e7134a_;
assign bus_00c9542f_=and_00b20115_u0;
assign or_00278af0_u0=bus_01ab54eb_|done_qual_u60_u0;
assign or_019749b6_u0=bus_01ab54eb_|bus_0144f414_|bus_01a25756_;
assign not_003da544_u0=~bus_0046cd71_;
assign mux_00427167_u0=({32{bus_01ab54eb_}}&bus_00eeb7ef_)|({32{bus_0144f414_}}&bus_00fee334_)|({32{bus_01a25756_}}&bus_003ad8b6_);
assign not_0149a6f6_u0=~bus_0046cd71_;
assign or_008914da_u0=bus_01ab54eb_|bus_0144f414_;
endmodule



module PROCESS_scheduler(CLK, RESET, GO, port_0182596d_, port_0148d67c_, port_015a802e_, port_01ead277_, port_00082475_, port_0041cb2b_, port_00795ad5_, port_01ac2e8e_, port_0059f665_, port_01c6ea35_, port_017d6741_, port_008097c7_, port_012cd222_, port_0195d97b_, RESULT, RESULT_u975, RESULT_u976, RESULT_u977, RESULT_u978, RESULT_u979, RESULT_u980, RESULT_u981, RESULT_u982, RESULT_u983, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_0182596d_;
input		port_0148d67c_;
input		port_015a802e_;
input	[31:0]	port_01ead277_;
input		port_00082475_;
input		port_0041cb2b_;
input		port_00795ad5_;
input		port_01ac2e8e_;
input		port_0059f665_;
input		port_01c6ea35_;
input		port_017d6741_;
input		port_008097c7_;
input		port_012cd222_;
input		port_0195d97b_;
output		RESULT;
output		RESULT_u975;
output		RESULT_u976;
output		RESULT_u977;
output		RESULT_u978;
output		RESULT_u979;
output		RESULT_u980;
output		RESULT_u981;
output		RESULT_u982;
output		RESULT_u983;
output		DONE;
wire		and_u1410_u0;
wire		and_u1411_u0;
wire		equals;
wire signed	[31:0]	equals_b_signed;
wire signed	[31:0]	equals_a_signed;
wire		and_u1412_u0;
wire		and_u1413_u0;
wire		and_u1414_u0;
wire		and_u1415_u0;
wire		not_u314_u0;
wire		not_u315_u0;
wire		and_u1416_u0;
wire		and_u1417_u0;
wire		simplePinWrite;
wire		and_u1418_u0;
wire		not_u316_u0;
wire		and_u1419_u0;
wire		and_u1420_u0;
wire		simplePinWrite_u418;
wire		and_u1421_u0;
reg		reg_0012a671_u0=1'h0;
reg		reg_01cdda0b_u0=1'h0;
wire		and_u1422_u0;
reg		reg_00f02141_u0=1'h0;
wire		or_u329_u0;
wire		and_u1423_u0;
wire		or_u330_u0;
wire		and_u1424_u0;
wire		and_u1425_u0;
reg		and_delayed_u24=1'h0;
wire		and_u1426_u0;
reg		and_delayed_u25_u0=1'h0;
wire		and_u1427_u0;
wire		or_u331_u0;
wire		and_u1428_u0;
wire		and_u1429_u0;
wire		not_u317_u0;
wire		simplePinWrite_u419;
wire		and_u1430_u0;
wire		and_u1431_u0;
wire		or_u332_u0;
wire		and_u1432_u0;
reg		reg_011995ce_u0=1'h0;
wire		and_u1433_u0;
wire		not_u318_u0;
wire		and_u1434_u0;
wire		and_u1435_u0;
wire		and_u1436_u0;
wire		and_u1437_u0;
wire		not_u319_u0;
wire		simplePinWrite_u420;
wire		and_u1438_u0;
wire		not_u320_u0;
wire		and_u1439_u0;
wire		and_u1440_u0;
wire		simplePinWrite_u421;
wire		and_u1441_u0;
reg		reg_01c8331d_u0=1'h0;
wire		or_u333_u0;
reg		and_delayed_u26_u0=1'h0;
reg		reg_0175ff81_u0=1'h0;
wire		and_u1442_u0;
wire		and_u1443_u0;
reg		reg_0135e90e_u0=1'h0;
wire		and_u1444_u0;
wire		or_u334_u0;
wire		and_u1445_u0;
reg		reg_00ac07fa_u0=1'h0;
wire		or_u335_u0;
wire		and_u1446_u0;
wire		and_u1447_u0;
wire		bus_018849a9_;
wire		scoreboard_01d9c592_resOr0;
wire		scoreboard_01d9c592_and;
wire		scoreboard_01d9c592_resOr1;
reg		scoreboard_01d9c592_reg2=1'h0;
reg		scoreboard_01d9c592_reg1=1'h0;
reg		scoreboard_01d9c592_reg0=1'h0;
wire		scoreboard_01d9c592_resOr2;
wire		or_u336_u0;
wire		mux_u248;
wire		doneCountIm_go_merge;
wire		or_u337_u0;
wire		mux_u249_u0;
wire		mux_u250_u0;
wire		or_u338_u0;
reg		syncEnable_u132=1'h0;
reg		syncEnable_u133_u0=1'h0;
reg		syncEnable_u134_u0=1'h0;
reg		syncEnable_u135_u0=1'h0;
reg		syncEnable_u136_u0=1'h0;
reg		block_GO_delayed_u14=1'h0;
wire		and_u1448_u0;
wire		or_u339_u0;
wire		or_u340_u0;
wire		mux_u251_u0;
reg		reg_01618569_u0=1'h0;
reg		reg_01618569_result_delayed_u0=1'h0;
wire		or_u341_u0;
wire		mux_u252_u0;
wire		mux_u253_u0;
wire		or_u342_u0;
assign and_u1410_u0=port_00795ad5_&port_012cd222_;
assign and_u1411_u0=and_u1410_u0&port_00082475_;
assign equals_a_signed=port_01ead277_;
assign equals_b_signed=32'h90;
assign equals=equals_a_signed==equals_b_signed;
assign and_u1412_u0=port_017d6741_&port_008097c7_;
assign and_u1413_u0=and_u1412_u0&port_0041cb2b_;
assign and_u1414_u0=block_GO_delayed_u14&not_u314_u0;
assign and_u1415_u0=block_GO_delayed_u14&syncEnable_u133_u0;
assign not_u314_u0=~syncEnable_u133_u0;
assign not_u315_u0=~syncEnable_u136_u0;
assign and_u1416_u0=and_u1427_u0&not_u315_u0;
assign and_u1417_u0=and_u1427_u0&syncEnable_u136_u0;
assign simplePinWrite=and_u1418_u0&{1{and_u1418_u0}};
assign and_u1418_u0=and_u1424_u0&and_u1424_u0;
assign not_u316_u0=~syncEnable_u132;
assign and_u1419_u0=and_u1425_u0&not_u316_u0;
assign and_u1420_u0=and_u1425_u0&syncEnable_u132;
assign simplePinWrite_u418=and_u1421_u0&{1{and_u1421_u0}};
assign and_u1421_u0=and_u1422_u0&and_u1422_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0012a671_u0<=1'h0;
else reg_0012a671_u0<=reg_01cdda0b_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01cdda0b_u0<=1'h0;
else reg_01cdda0b_u0<=and_u1422_u0;
end
assign and_u1422_u0=and_u1420_u0&and_u1425_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00f02141_u0<=1'h0;
else reg_00f02141_u0<=and_u1423_u0;
end
assign or_u329_u0=reg_00f02141_u0|reg_0012a671_u0;
assign and_u1423_u0=and_u1419_u0&and_u1425_u0;
assign or_u330_u0=and_delayed_u24|or_u329_u0;
assign and_u1424_u0=and_u1417_u0&and_u1427_u0;
assign and_u1425_u0=and_u1416_u0&and_u1427_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u24<=1'h0;
else and_delayed_u24<=and_u1424_u0;
end
assign and_u1426_u0=and_u1414_u0&block_GO_delayed_u14;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u25_u0<=1'h0;
else and_delayed_u25_u0<=and_u1426_u0;
end
assign and_u1427_u0=and_u1415_u0&block_GO_delayed_u14;
assign or_u331_u0=or_u330_u0|and_delayed_u25_u0;
assign and_u1428_u0=block_GO_delayed_u14&not_u317_u0;
assign and_u1429_u0=block_GO_delayed_u14&syncEnable_u135_u0;
assign not_u317_u0=~syncEnable_u135_u0;
assign simplePinWrite_u419=and_u1430_u0&{1{and_u1430_u0}};
assign and_u1430_u0=and_u1431_u0&and_u1431_u0;
assign and_u1431_u0=and_u1432_u0&and_u1432_u0;
assign or_u332_u0=reg_011995ce_u0|port_0195d97b_;
assign and_u1432_u0=and_u1429_u0&block_GO_delayed_u14;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_011995ce_u0<=1'h0;
else reg_011995ce_u0<=and_u1433_u0;
end
assign and_u1433_u0=and_u1428_u0&block_GO_delayed_u14;
assign not_u318_u0=~syncEnable_u134_u0;
assign and_u1434_u0=block_GO_delayed_u14&not_u318_u0;
assign and_u1435_u0=block_GO_delayed_u14&syncEnable_u134_u0;
assign and_u1436_u0=and_u1447_u0&syncEnable_u136_u0;
assign and_u1437_u0=and_u1447_u0&not_u319_u0;
assign not_u319_u0=~syncEnable_u136_u0;
assign simplePinWrite_u420=and_u1438_u0&{1{and_u1438_u0}};
assign and_u1438_u0=and_u1445_u0&and_u1445_u0;
assign not_u320_u0=~and_u1413_u0;
assign and_u1439_u0=and_u1443_u0&and_u1413_u0;
assign and_u1440_u0=and_u1443_u0&not_u320_u0;
assign simplePinWrite_u421=and_u1442_u0&{1{and_u1442_u0}};
assign and_u1441_u0=and_u1440_u0&and_u1443_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01c8331d_u0<=1'h0;
else reg_01c8331d_u0<=reg_0175ff81_u0;
end
assign or_u333_u0=and_delayed_u26_u0|reg_01c8331d_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u26_u0<=1'h0;
else and_delayed_u26_u0<=and_u1441_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0175ff81_u0<=1'h0;
else reg_0175ff81_u0<=and_u1442_u0;
end
assign and_u1442_u0=and_u1439_u0&and_u1443_u0;
assign and_u1443_u0=and_u1444_u0&and_u1444_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0135e90e_u0<=1'h0;
else reg_0135e90e_u0<=and_u1445_u0;
end
assign and_u1444_u0=and_u1437_u0&and_u1447_u0;
assign or_u334_u0=or_u333_u0|reg_0135e90e_u0;
assign and_u1445_u0=and_u1436_u0&and_u1447_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00ac07fa_u0<=1'h0;
else reg_00ac07fa_u0<=and_u1446_u0;
end
assign or_u335_u0=reg_00ac07fa_u0|or_u334_u0;
assign and_u1446_u0=and_u1434_u0&block_GO_delayed_u14;
assign and_u1447_u0=and_u1435_u0&block_GO_delayed_u14;
assign bus_018849a9_=scoreboard_01d9c592_and|RESET;
assign scoreboard_01d9c592_resOr0=or_u331_u0|scoreboard_01d9c592_reg0;
assign scoreboard_01d9c592_and=scoreboard_01d9c592_resOr0&scoreboard_01d9c592_resOr1&scoreboard_01d9c592_resOr2;
assign scoreboard_01d9c592_resOr1=or_u332_u0|scoreboard_01d9c592_reg1;
always @(posedge CLK)
begin
if (bus_018849a9_)
scoreboard_01d9c592_reg2<=1'h0;
else if (or_u335_u0)
scoreboard_01d9c592_reg2<=1'h1;
else scoreboard_01d9c592_reg2<=scoreboard_01d9c592_reg2;
end
always @(posedge CLK)
begin
if (bus_018849a9_)
scoreboard_01d9c592_reg1<=1'h0;
else if (or_u332_u0)
scoreboard_01d9c592_reg1<=1'h1;
else scoreboard_01d9c592_reg1<=scoreboard_01d9c592_reg1;
end
always @(posedge CLK)
begin
if (bus_018849a9_)
scoreboard_01d9c592_reg0<=1'h0;
else if (or_u331_u0)
scoreboard_01d9c592_reg0<=1'h1;
else scoreboard_01d9c592_reg0<=scoreboard_01d9c592_reg0;
end
assign scoreboard_01d9c592_resOr2=or_u335_u0|scoreboard_01d9c592_reg2;
assign or_u336_u0=and_u1430_u0|and_u1438_u0;
assign mux_u248=(and_u1430_u0)?1'h1:1'h0;
assign doneCountIm_go_merge=simplePinWrite|simplePinWrite_u420;
assign or_u337_u0=and_u1418_u0|and_u1430_u0;
assign mux_u249_u0=(and_u1418_u0)?1'h1:1'h0;
assign mux_u250_u0=(and_u1418_u0)?1'h0:1'h1;
assign or_u338_u0=and_u1418_u0|and_u1438_u0;
always @(posedge CLK)
begin
if (and_u1448_u0)
syncEnable_u132<=and_u1411_u0;
end
always @(posedge CLK)
begin
if (and_u1448_u0)
syncEnable_u133_u0<=port_0182596d_;
end
always @(posedge CLK)
begin
if (and_u1448_u0)
syncEnable_u134_u0<=port_015a802e_;
end
always @(posedge CLK)
begin
if (and_u1448_u0)
syncEnable_u135_u0<=port_0148d67c_;
end
always @(posedge CLK)
begin
if (and_u1448_u0)
syncEnable_u136_u0<=equals;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u14<=1'h0;
else block_GO_delayed_u14<=and_u1448_u0;
end
assign and_u1448_u0=or_u339_u0&or_u339_u0;
assign or_u339_u0=reg_01618569_result_delayed_u0|scoreboard_01d9c592_and;
assign or_u340_u0=GO|or_u336_u0;
assign mux_u251_u0=(GO)?1'h0:mux_u248;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01618569_u0<=1'h0;
else reg_01618569_u0<=GO;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01618569_result_delayed_u0<=1'h0;
else reg_01618569_result_delayed_u0<=reg_01618569_u0;
end
assign or_u341_u0=GO|or_u338_u0;
assign mux_u252_u0=(GO)?1'h1:mux_u250_u0;
assign mux_u253_u0=(GO)?1'h0:mux_u249_u0;
assign or_u342_u0=GO|or_u337_u0;
assign RESULT=or_u341_u0;
assign RESULT_u975=mux_u252_u0;
assign RESULT_u976=or_u342_u0;
assign RESULT_u977=mux_u253_u0;
assign RESULT_u978=or_u340_u0;
assign RESULT_u979=mux_u251_u0;
assign RESULT_u980=simplePinWrite_u421;
assign RESULT_u981=simplePinWrite_u419;
assign RESULT_u982=doneCountIm_go_merge;
assign RESULT_u983=simplePinWrite_u418;
assign DONE=1'h0;
endmodule



module PROCESS_structuralmemory_00814577_(CLK_u17, bus_01c52148_, bus_00890cb8_, bus_014efb86_, bus_00aef9ca_, bus_00e5479e_, bus_010d9e31_, bus_0000f23b_, bus_00b89a1d_, bus_01d3fa4a_, bus_0118cc44_, bus_019151a3_, bus_010cc662_, bus_010aabe7_);
input		CLK_u17;
input		bus_01c52148_;
input	[31:0]	bus_00890cb8_;
input	[2:0]	bus_014efb86_;
input		bus_00aef9ca_;
input		bus_00e5479e_;
input	[7:0]	bus_010d9e31_;
input	[31:0]	bus_0000f23b_;
input	[2:0]	bus_00b89a1d_;
input		bus_01d3fa4a_;
input	[7:0]	bus_0118cc44_;
output	[7:0]	bus_019151a3_;
output		bus_010cc662_;
output		bus_010aabe7_;
wire		or_01ae1400_u0;
reg		logicalMem_38cddc_we_delay0_u0=1'h0;
reg		logicalMem_38cddc_re_delay0_u0=1'h0;
wire	[7:0]	bus_01900bb9_;
reg		logicalMem_38cddc_we_delay0_u1_u0=1'h0;
wire		or_00f88af3_u0;
assign or_01ae1400_u0=logicalMem_38cddc_re_delay0_u0|logicalMem_38cddc_we_delay0_u0;
always @(posedge CLK_u17 or posedge bus_01c52148_)
begin
if (bus_01c52148_)
logicalMem_38cddc_we_delay0_u0<=1'h0;
else logicalMem_38cddc_we_delay0_u0<=bus_00e5479e_;
end
always @(posedge CLK_u17 or posedge bus_01c52148_)
begin
if (bus_01c52148_)
logicalMem_38cddc_re_delay0_u0<=1'h0;
else logicalMem_38cddc_re_delay0_u0<=bus_00aef9ca_;
end
assign bus_019151a3_=bus_01900bb9_;
assign bus_010cc662_=or_01ae1400_u0;
assign bus_010aabe7_=logicalMem_38cddc_we_delay0_u1_u0;
PROCESS_forge_memory_25344x8_27 PROCESS_forge_memory_25344x8_27_instance1(.CLK(CLK_u17), 
  .ENA(or_00f88af3_u0), .WEA(bus_00e5479e_), .DINA(bus_010d9e31_), .ADDRA(bus_00890cb8_), 
  .DOUTA(bus_01900bb9_), .DONEA(), .ENB(bus_01d3fa4a_), .WEB(bus_01d3fa4a_), .DINB(8'h0), 
  .ADDRB(bus_0000f23b_), .DONEB());
always @(posedge CLK_u17 or posedge bus_01c52148_)
begin
if (bus_01c52148_)
logicalMem_38cddc_we_delay0_u1_u0<=1'h0;
else logicalMem_38cddc_we_delay0_u1_u0<=bus_01d3fa4a_;
end
assign or_00f88af3_u0=bus_00aef9ca_|bus_00e5479e_;
endmodule



module PROCESS_drawRectangle(CLK, RESET, GO, port_0130bfa1_, port_01243a78_, port_006015e8_, port_014d58fd_, port_01cb501c_, port_00e850d8_, RESULT, RESULT_u984, RESULT_u985, RESULT_u986, RESULT_u987, RESULT_u988, RESULT_u989, RESULT_u990, RESULT_u991, RESULT_u992, RESULT_u993, RESULT_u994, RESULT_u995, RESULT_u996, RESULT_u997, RESULT_u998, RESULT_u999, RESULT_u1000, RESULT_u1001, RESULT_u1002, RESULT_u1003, RESULT_u1004, RESULT_u1005, RESULT_u1006, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_0130bfa1_;
input		port_01243a78_;
input		port_006015e8_;
input		port_014d58fd_;
input		port_01cb501c_;
input		port_00e850d8_;
output		RESULT;
output	[31:0]	RESULT_u984;
output	[7:0]	RESULT_u985;
output	[2:0]	RESULT_u986;
output		RESULT_u987;
output	[31:0]	RESULT_u988;
output	[7:0]	RESULT_u989;
output	[2:0]	RESULT_u990;
output		RESULT_u991;
output	[31:0]	RESULT_u992;
output	[7:0]	RESULT_u993;
output	[2:0]	RESULT_u994;
output		RESULT_u995;
output	[31:0]	RESULT_u996;
output	[7:0]	RESULT_u997;
output	[2:0]	RESULT_u998;
output		RESULT_u999;
output	[31:0]	RESULT_u1000;
output	[7:0]	RESULT_u1001;
output	[2:0]	RESULT_u1002;
output		RESULT_u1003;
output	[31:0]	RESULT_u1004;
output	[7:0]	RESULT_u1005;
output	[2:0]	RESULT_u1006;
output		DONE;
reg		reg_009197a7_u0=1'h0;
wire	[31:0]	add;
wire	[31:0]	add_u524;
reg		reg_00323d5a_u0=1'h0;
wire		or_u343_u0;
wire		and_u1449_u0;
wire	[31:0]	add_u525;
wire	[31:0]	add_u526;
wire		or_u344_u0;
wire		and_u1450_u0;
reg		reg_008228c8_u0=1'h0;
wire	[31:0]	add_u527;
wire	[31:0]	add_u528;
reg		reg_007ed15f_u0=1'h0;
wire		or_u345_u0;
wire		and_u1451_u0;
wire	[31:0]	add_u529;
wire	[31:0]	add_u530;
wire		or_u346_u0;
reg		reg_01648375_u0=1'h0;
wire		and_u1452_u0;
wire	[31:0]	add_u531;
wire	[31:0]	add_u532;
reg		reg_00b62503_u0=1'h0;
wire		and_u1453_u0;
wire		or_u347_u0;
wire	[31:0]	add_u533;
wire	[31:0]	add_u534;
wire		or_u348_u0;
reg		reg_00f560a5_u0=1'h0;
wire		and_u1454_u0;
wire	[31:0]	add_u535;
reg	[31:0]	syncEnable_u137=32'h0;
reg	[31:0]	syncEnable_u138_u0=32'h0;
reg	[31:0]	syncEnable_u139_u0=32'h0;
reg	[31:0]	syncEnable_u140_u0=32'h0;
reg	[31:0]	syncEnable_u141_u0=32'h0;
reg	[31:0]	syncEnable_u142_u0=32'h0;
reg		block_GO_delayed_u15=1'h0;
reg		block_GO_delayed_result_delayed_u3=1'h0;
reg	[31:0]	syncEnable_u143_u0=32'h0;
wire		and_u1455_u0;
reg		reg_009197a7_result_delayed_u0=1'h0;
wire		lessThanEqualTo;
wire signed	[31:0]	lessThanEqualTo_b_signed;
wire signed	[31:0]	lessThanEqualTo_a_signed;
wire		and_u1456_u0;
wire		and_u1457_u0;
wire		not_u321_u0;
reg		reg_009197a7_result_delayed_result_delayed_u0=1'h0;
wire		and_u1458_u0;
wire	[31:0]	latch_0079af26_out;
reg	[6:0]	latch_0079af26_reg=7'h0;
wire		or_u349_u0;
wire	[31:0]	mux_u254;
wire		and_u1459_u0;
reg		and_delayed_u27=1'h0;
wire		and_u1460_u0;
wire	[31:0]	add_u536;
wire	[31:0]	add_u537;
wire	[31:0]	add_u538;
wire	[31:0]	add_u539;
reg		reg_01920b86_u0=1'h0;
wire		and_u1461_u0;
wire		or_u350_u0;
wire	[31:0]	add_u540;
wire	[31:0]	add_u541;
wire	[31:0]	add_u542;
wire	[31:0]	add_u543;
wire		or_u351_u0;
wire		and_u1462_u0;
reg		reg_00960b3f_u0=1'h0;
wire	[31:0]	add_u544;
wire	[31:0]	add_u545;
wire	[31:0]	add_u546;
wire	[31:0]	add_u547;
reg		reg_00f58588_u0=1'h0;
wire		or_u352_u0;
wire		and_u1463_u0;
wire	[31:0]	add_u548;
wire	[31:0]	add_u549;
wire	[31:0]	add_u550;
wire	[31:0]	add_u551;
wire		or_u353_u0;
wire		and_u1464_u0;
reg		reg_01e60b91_u0=1'h0;
wire	[31:0]	add_u552;
wire	[31:0]	add_u553;
wire	[31:0]	add_u554;
wire	[31:0]	add_u555;
wire		or_u354_u0;
wire		and_u1465_u0;
reg		reg_00af90bc_u0=1'h0;
wire	[31:0]	add_u556;
wire	[31:0]	add_u557;
wire	[31:0]	add_u558;
wire	[31:0]	add_u559;
wire		and_u1466_u0;
reg		reg_01b1224d_u0=1'h0;
wire		or_u355_u0;
wire	[31:0]	add_u560;
reg	[31:0]	syncEnable_u144_u0=32'h0;
reg	[31:0]	syncEnable_u145_u0=32'h0;
reg	[31:0]	syncEnable_u146_u0=32'h0;
reg	[31:0]	syncEnable_u147_u0=32'h0;
reg	[31:0]	syncEnable_u148_u0=32'h0;
reg	[31:0]	syncEnable_u149_u0=32'h0;
reg		reg_01c542a1_u0=1'h0;
reg	[31:0]	syncEnable_u150_u0=32'h0;
reg		block_GO_delayed_u16_u0=1'h0;
reg		reg_004c46af_u0=1'h0;
wire signed	[31:0]	lessThanEqualTo_u4_b_signed;
wire		lessThanEqualTo_u4;
wire signed	[31:0]	lessThanEqualTo_u4_a_signed;
wire		not_u322_u0;
wire		and_u1467_u0;
wire		and_u1468_u0;
reg		and_delayed_result_delayed_u2=1'h0;
wire		or_u356_u0;
wire	[31:0]	latch_009252a5_out;
reg	[6:0]	latch_009252a5_reg=7'h0;
wire	[31:0]	mux_u255_u0;
wire	[31:0]	latch_009976f9_out;
reg	[5:0]	latch_009976f9_reg=6'h0;
reg	[6:0]	latch_0113a81c_reg=7'h0;
wire	[31:0]	latch_0113a81c_out;
wire		or_u357_u0;
wire	[31:0]	mux_u256_u0;
reg		reg_01b7cb8c_u0=1'h0;
wire		or_u358_u0;
wire	[31:0]	mux_u257_u0;
wire	[31:0]	mux_u258_u0;
wire		or_u359_u0;
wire		or_u360_u0;
wire	[31:0]	mux_u259_u0;
wire		or_u361_u0;
wire	[31:0]	mux_u260_u0;
wire	[31:0]	mux_u261_u0;
wire		or_u362_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_009197a7_u0<=1'h0;
else reg_009197a7_u0<=and_u1458_u0;
end
assign add=32'h1130+mux_u254;
assign add_u524=32'h0+add;
always @(posedge CLK or posedge block_GO_delayed_u15 or posedge or_u343_u0)
begin
if (or_u343_u0)
reg_00323d5a_u0<=1'h0;
else if (block_GO_delayed_u15)
reg_00323d5a_u0<=1'h1;
else reg_00323d5a_u0<=reg_00323d5a_u0;
end
assign or_u343_u0=and_u1449_u0|RESET;
assign and_u1449_u0=reg_00323d5a_u0&port_006015e8_;
assign add_u525=32'h1130+mux_u254;
assign add_u526=32'h0+add_u525;
assign or_u344_u0=and_u1450_u0|RESET;
assign and_u1450_u0=reg_008228c8_u0&port_01243a78_;
always @(posedge CLK or posedge block_GO_delayed_u15 or posedge or_u344_u0)
begin
if (or_u344_u0)
reg_008228c8_u0<=1'h0;
else if (block_GO_delayed_u15)
reg_008228c8_u0<=1'h1;
else reg_008228c8_u0<=reg_008228c8_u0;
end
assign add_u527=32'h1130+mux_u254;
assign add_u528=32'h0+add_u527;
always @(posedge CLK or posedge block_GO_delayed_u15 or posedge or_u345_u0)
begin
if (or_u345_u0)
reg_007ed15f_u0<=1'h0;
else if (block_GO_delayed_u15)
reg_007ed15f_u0<=1'h1;
else reg_007ed15f_u0<=reg_007ed15f_u0;
end
assign or_u345_u0=and_u1451_u0|RESET;
assign and_u1451_u0=reg_007ed15f_u0&port_0130bfa1_;
assign add_u529=32'h25d0+mux_u254;
assign add_u530=32'h0+add_u529;
assign or_u346_u0=and_u1452_u0|RESET;
always @(posedge CLK or posedge block_GO_delayed_result_delayed_u3 or posedge or_u346_u0)
begin
if (or_u346_u0)
reg_01648375_u0<=1'h0;
else if (block_GO_delayed_result_delayed_u3)
reg_01648375_u0<=1'h1;
else reg_01648375_u0<=reg_01648375_u0;
end
assign and_u1452_u0=reg_01648375_u0&port_01cb501c_;
assign add_u531=32'h25d0+mux_u254;
assign add_u532=32'h0+add_u531;
always @(posedge CLK or posedge block_GO_delayed_result_delayed_u3 or posedge or_u347_u0)
begin
if (or_u347_u0)
reg_00b62503_u0<=1'h0;
else if (block_GO_delayed_result_delayed_u3)
reg_00b62503_u0<=1'h1;
else reg_00b62503_u0<=reg_00b62503_u0;
end
assign and_u1453_u0=reg_00b62503_u0&port_014d58fd_;
assign or_u347_u0=and_u1453_u0|RESET;
assign add_u533=32'h25d0+mux_u254;
assign add_u534=32'h0+add_u533;
assign or_u348_u0=and_u1454_u0|RESET;
always @(posedge CLK or posedge block_GO_delayed_result_delayed_u3 or posedge or_u348_u0)
begin
if (or_u348_u0)
reg_00f560a5_u0<=1'h0;
else if (block_GO_delayed_result_delayed_u3)
reg_00f560a5_u0<=1'h1;
else reg_00f560a5_u0<=reg_00f560a5_u0;
end
assign and_u1454_u0=reg_00f560a5_u0&port_00e850d8_;
assign add_u535=mux_u254+32'h1;
always @(posedge CLK)
begin
if (and_u1458_u0)
syncEnable_u137<=add_u528;
end
always @(posedge CLK)
begin
if (and_u1458_u0)
syncEnable_u138_u0<=add_u530;
end
always @(posedge CLK)
begin
if (and_u1458_u0)
syncEnable_u139_u0<=add_u524;
end
always @(posedge CLK)
begin
if (and_u1458_u0)
syncEnable_u140_u0<=add_u526;
end
always @(posedge CLK)
begin
if (and_u1458_u0)
syncEnable_u141_u0<=add_u534;
end
always @(posedge CLK)
begin
if (and_u1458_u0)
syncEnable_u142_u0<=add_u532;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u15<=1'h0;
else block_GO_delayed_u15<=and_u1458_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_result_delayed_u3<=1'h0;
else block_GO_delayed_result_delayed_u3<=block_GO_delayed_u15;
end
always @(posedge CLK)
begin
if (and_u1458_u0)
syncEnable_u143_u0<=add_u535;
end
assign and_u1455_u0=and_u1457_u0&or_u349_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_009197a7_result_delayed_u0<=1'h0;
else reg_009197a7_result_delayed_u0<=reg_009197a7_u0;
end
assign lessThanEqualTo_a_signed=mux_u254;
assign lessThanEqualTo_b_signed=32'h32;
assign lessThanEqualTo=lessThanEqualTo_a_signed<=lessThanEqualTo_b_signed;
assign and_u1456_u0=or_u349_u0&lessThanEqualTo;
assign and_u1457_u0=or_u349_u0&not_u321_u0;
assign not_u321_u0=~lessThanEqualTo;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_009197a7_result_delayed_result_delayed_u0<=1'h0;
else reg_009197a7_result_delayed_result_delayed_u0<=reg_009197a7_result_delayed_u0;
end
assign and_u1458_u0=and_u1456_u0&or_u349_u0;
assign latch_0079af26_out=(reg_01b7cb8c_u0)?32'h32:32'h32;
always @(posedge CLK)
begin
if (reg_01b7cb8c_u0)
latch_0079af26_reg<=7'h32;
end
assign or_u349_u0=reg_009197a7_result_delayed_result_delayed_u0|reg_01b7cb8c_u0;
assign mux_u254=(reg_009197a7_result_delayed_result_delayed_u0)?syncEnable_u143_u0:32'h1e;
assign and_u1459_u0=and_u1468_u0&or_u356_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u27<=1'h0;
else and_delayed_u27<=and_u1459_u0;
end
assign and_u1460_u0=and_u1467_u0&or_u356_u0;
assign add_u536={mux_u255_u0[24:0], 7'b0}+{mux_u255_u0[26:0], 5'b0};
assign add_u537={add_u536[31:5], 5'b0}+{mux_u255_u0[27:0], 4'b0};
assign add_u538={add_u537[31:4], 4'b0}+32'h1e;
assign add_u539=32'h0+{add_u538[31:4], 4'b1110};
always @(posedge CLK or posedge block_GO_delayed_u16_u0 or posedge or_u350_u0)
begin
if (or_u350_u0)
reg_01920b86_u0<=1'h0;
else if (block_GO_delayed_u16_u0)
reg_01920b86_u0<=1'h1;
else reg_01920b86_u0<=reg_01920b86_u0;
end
assign and_u1461_u0=reg_01920b86_u0&port_006015e8_;
assign or_u350_u0=and_u1461_u0|RESET;
assign add_u540={mux_u255_u0[24:0], 7'b0}+{mux_u255_u0[26:0], 5'b0};
assign add_u541={add_u540[31:5], 5'b0}+{mux_u255_u0[27:0], 4'b0};
assign add_u542={add_u541[31:4], 4'b0}+32'h1e;
assign add_u543=32'h0+{add_u542[31:4], 4'b1110};
assign or_u351_u0=and_u1462_u0|RESET;
assign and_u1462_u0=reg_00960b3f_u0&port_01243a78_;
always @(posedge CLK or posedge block_GO_delayed_u16_u0 or posedge or_u351_u0)
begin
if (or_u351_u0)
reg_00960b3f_u0<=1'h0;
else if (block_GO_delayed_u16_u0)
reg_00960b3f_u0<=1'h1;
else reg_00960b3f_u0<=reg_00960b3f_u0;
end
assign add_u544={mux_u255_u0[24:0], 7'b0}+{mux_u255_u0[26:0], 5'b0};
assign add_u545={add_u544[31:5], 5'b0}+{mux_u255_u0[27:0], 4'b0};
assign add_u546={add_u545[31:4], 4'b0}+32'h1e;
assign add_u547=32'h0+{add_u546[31:4], 4'b1110};
always @(posedge CLK or posedge block_GO_delayed_u16_u0 or posedge or_u352_u0)
begin
if (or_u352_u0)
reg_00f58588_u0<=1'h0;
else if (block_GO_delayed_u16_u0)
reg_00f58588_u0<=1'h1;
else reg_00f58588_u0<=reg_00f58588_u0;
end
assign or_u352_u0=and_u1463_u0|RESET;
assign and_u1463_u0=reg_00f58588_u0&port_0130bfa1_;
assign add_u548={mux_u255_u0[24:0], 7'b0}+{mux_u255_u0[26:0], 5'b0};
assign add_u549={add_u548[31:5], 5'b0}+{mux_u255_u0[27:0], 4'b0};
assign add_u550={add_u549[31:4], 4'b0}+32'h32;
assign add_u551=32'h0+{add_u550[31:4], 4'b10};
assign or_u353_u0=and_u1464_u0|RESET;
assign and_u1464_u0=reg_01e60b91_u0&port_01cb501c_;
always @(posedge CLK or posedge reg_01c542a1_u0 or posedge or_u353_u0)
begin
if (or_u353_u0)
reg_01e60b91_u0<=1'h0;
else if (reg_01c542a1_u0)
reg_01e60b91_u0<=1'h1;
else reg_01e60b91_u0<=reg_01e60b91_u0;
end
assign add_u552={mux_u255_u0[24:0], 7'b0}+{mux_u255_u0[26:0], 5'b0};
assign add_u553={add_u552[31:5], 5'b0}+{mux_u255_u0[27:0], 4'b0};
assign add_u554={add_u553[31:4], 4'b0}+32'h32;
assign add_u555=32'h0+{add_u554[31:4], 4'b10};
assign or_u354_u0=and_u1465_u0|RESET;
assign and_u1465_u0=reg_00af90bc_u0&port_014d58fd_;
always @(posedge CLK or posedge reg_01c542a1_u0 or posedge or_u354_u0)
begin
if (or_u354_u0)
reg_00af90bc_u0<=1'h0;
else if (reg_01c542a1_u0)
reg_00af90bc_u0<=1'h1;
else reg_00af90bc_u0<=reg_00af90bc_u0;
end
assign add_u556={mux_u255_u0[24:0], 7'b0}+{mux_u255_u0[26:0], 5'b0};
assign add_u557={add_u556[31:5], 5'b0}+{mux_u255_u0[27:0], 4'b0};
assign add_u558={add_u557[31:4], 4'b0}+32'h32;
assign add_u559=32'h0+{add_u558[31:4], 4'b10};
assign and_u1466_u0=reg_01b1224d_u0&port_00e850d8_;
always @(posedge CLK or posedge reg_01c542a1_u0 or posedge or_u355_u0)
begin
if (or_u355_u0)
reg_01b1224d_u0<=1'h0;
else if (reg_01c542a1_u0)
reg_01b1224d_u0<=1'h1;
else reg_01b1224d_u0<=reg_01b1224d_u0;
end
assign or_u355_u0=and_u1466_u0|RESET;
assign add_u560=mux_u255_u0+32'h1;
always @(posedge CLK)
begin
if (and_u1459_u0)
syncEnable_u144_u0<={add_u547[31:4], 4'b1110};
end
always @(posedge CLK)
begin
if (and_u1459_u0)
syncEnable_u145_u0<={add_u559[31:4], 4'b10};
end
always @(posedge CLK)
begin
if (and_u1459_u0)
syncEnable_u146_u0<={add_u539[31:4], 4'b1110};
end
always @(posedge CLK)
begin
if (and_u1459_u0)
syncEnable_u147_u0<={add_u551[31:4], 4'b10};
end
always @(posedge CLK)
begin
if (and_u1459_u0)
syncEnable_u148_u0<={add_u543[31:4], 4'b1110};
end
always @(posedge CLK)
begin
if (and_u1459_u0)
syncEnable_u149_u0<=add_u560;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01c542a1_u0<=1'h0;
else reg_01c542a1_u0<=block_GO_delayed_u16_u0;
end
always @(posedge CLK)
begin
if (and_u1459_u0)
syncEnable_u150_u0<={add_u555[31:4], 4'b10};
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u16_u0<=1'h0;
else block_GO_delayed_u16_u0<=and_u1459_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_004c46af_u0<=1'h0;
else reg_004c46af_u0<=and_delayed_result_delayed_u2;
end
assign lessThanEqualTo_u4_a_signed=mux_u255_u0;
assign lessThanEqualTo_u4_b_signed=32'h37;
assign lessThanEqualTo_u4=lessThanEqualTo_u4_a_signed<=lessThanEqualTo_u4_b_signed;
assign not_u322_u0=~lessThanEqualTo_u4;
assign and_u1467_u0=or_u356_u0&not_u322_u0;
assign and_u1468_u0=or_u356_u0&lessThanEqualTo_u4;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_result_delayed_u2<=1'h0;
else and_delayed_result_delayed_u2<=and_delayed_u27;
end
assign or_u356_u0=reg_004c46af_u0|and_u1455_u0;
assign latch_009252a5_out=(and_u1455_u0)?32'h37:32'h37;
always @(posedge CLK)
begin
if (and_u1455_u0)
latch_009252a5_reg<=7'h37;
end
assign mux_u255_u0=(reg_004c46af_u0)?syncEnable_u149_u0:32'h19;
assign latch_009976f9_out=(and_u1455_u0)?32'h1e:32'h1e;
always @(posedge CLK)
begin
if (and_u1455_u0)
latch_009976f9_reg<=6'h1e;
end
always @(posedge CLK)
begin
if (and_u1455_u0)
latch_0113a81c_reg<=7'h32;
end
assign latch_0113a81c_out=(and_u1455_u0)?32'h32:32'h32;
assign or_u357_u0=block_GO_delayed_result_delayed_u3|reg_01c542a1_u0;
assign mux_u256_u0=(block_GO_delayed_result_delayed_u3)?syncEnable_u138_u0:{syncEnable_u147_u0[31:4], 4'b10};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01b7cb8c_u0<=1'h0;
else reg_01b7cb8c_u0<=GO;
end
assign or_u358_u0=block_GO_delayed_result_delayed_u3|reg_01c542a1_u0;
assign mux_u257_u0=(block_GO_delayed_result_delayed_u3)?syncEnable_u142_u0:{syncEnable_u150_u0[31:4], 4'b10};
assign mux_u258_u0=(block_GO_delayed_u15)?syncEnable_u137:{syncEnable_u144_u0[31:4], 4'b1110};
assign or_u359_u0=block_GO_delayed_u15|block_GO_delayed_u16_u0;
assign or_u360_u0=block_GO_delayed_result_delayed_u3|reg_01c542a1_u0;
assign mux_u259_u0=(block_GO_delayed_result_delayed_u3)?syncEnable_u141_u0:{syncEnable_u145_u0[31:4], 4'b10};
assign or_u361_u0=block_GO_delayed_u15|block_GO_delayed_u16_u0;
assign mux_u260_u0=(block_GO_delayed_u15)?syncEnable_u140_u0:{syncEnable_u148_u0[31:4], 4'b1110};
assign mux_u261_u0=(block_GO_delayed_u15)?syncEnable_u139_u0:{syncEnable_u146_u0[31:4], 4'b1110};
assign or_u362_u0=block_GO_delayed_u15|block_GO_delayed_u16_u0;
assign RESULT=or_u359_u0;
assign RESULT_u984=mux_u258_u0;
assign RESULT_u985=8'h0;
assign RESULT_u986=3'h1;
assign RESULT_u987=or_u361_u0;
assign RESULT_u988=mux_u260_u0;
assign RESULT_u989=8'h0;
assign RESULT_u990=3'h1;
assign RESULT_u991=or_u362_u0;
assign RESULT_u992=mux_u261_u0;
assign RESULT_u993=8'hff;
assign RESULT_u994=3'h1;
assign RESULT_u995=or_u358_u0;
assign RESULT_u996=mux_u257_u0;
assign RESULT_u997=8'h0;
assign RESULT_u998=3'h1;
assign RESULT_u999=or_u357_u0;
assign RESULT_u1000=mux_u256_u0;
assign RESULT_u1001=8'hff;
assign RESULT_u1002=3'h1;
assign RESULT_u1003=or_u360_u0;
assign RESULT_u1004=mux_u259_u0;
assign RESULT_u1005=8'h0;
assign RESULT_u1006=3'h1;
assign DONE=and_u1460_u0;
endmodule



module PROCESS_send(CLK, RESET, GO, port_01245fcb_, port_00c7b822_, port_00817c5e_, port_015914f6_, port_010e3311_, port_0148441b_, port_012755fe_, port_0041b215_, RESULT, RESULT_u1007, RESULT_u1008, RESULT_u1009, RESULT_u1010, RESULT_u1011, RESULT_u1012, RESULT_u1013, RESULT_u1014, RESULT_u1015, RESULT_u1016, RESULT_u1017, RESULT_u1018, RESULT_u1019, RESULT_u1020, RESULT_u1021, RESULT_u1022, RESULT_u1023, RESULT_u1024, RESULT_u1025, RESULT_u1026, RESULT_u1027, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_01245fcb_;
input	[31:0]	port_00c7b822_;
input		port_00817c5e_;
input	[7:0]	port_015914f6_;
input		port_010e3311_;
input	[7:0]	port_0148441b_;
input		port_012755fe_;
input	[7:0]	port_0041b215_;
output		RESULT;
output	[31:0]	RESULT_u1007;
output		RESULT_u1008;
output	[31:0]	RESULT_u1009;
output		RESULT_u1010;
output	[31:0]	RESULT_u1011;
output	[2:0]	RESULT_u1012;
output		RESULT_u1013;
output	[31:0]	RESULT_u1014;
output	[2:0]	RESULT_u1015;
output		RESULT_u1016;
output	[31:0]	RESULT_u1017;
output	[2:0]	RESULT_u1018;
output	[7:0]	RESULT_u1019;
output	[15:0]	RESULT_u1020;
output	[15:0]	RESULT_u1021;
output	[7:0]	RESULT_u1022;
output		RESULT_u1023;
output		RESULT_u1024;
output		RESULT_u1025;
output	[15:0]	RESULT_u1026;
output	[7:0]	RESULT_u1027;
output		DONE;
wire	[31:0]	add;
wire	[31:0]	add_u561;
wire	[31:0]	add_u562;
wire	[31:0]	add_u563;
wire		or_u363_u0;
wire		and_u1469_u0;
reg		done_cache_u16=1'h0;
wire	[31:0]	add_u564;
wire	[31:0]	add_u565;
wire	[31:0]	add_u566;
wire	[31:0]	add_u567;
wire		or_u364_u0;
wire		and_u1470_u0;
reg		done_cache_u17_u0=1'h0;
wire	[31:0]	add_u568;
wire	[31:0]	add_u569;
wire	[31:0]	add_u570;
wire	[31:0]	add_u571;
wire		and_u1471_u0;
wire		or_u365_u0;
reg		done_cache_u18_u0=1'h0;
wire	[31:0]	add_u572;
wire signed	[31:0]	equals_a_signed;
wire signed	[31:0]	equals_b_signed;
wire		equals;
wire		and_u1472_u0;
wire		and_u1473_u0;
wire		not_u323_u0;
wire	[31:0]	add_u573;
wire	[31:0]	mux_u262;
wire		and_u1474_u0;
wire		and_u1475_u0;
wire	[31:0]	mux_u263_u0;
wire		simplePinWrite;
wire	[7:0]	simplePinWrite_u422;
wire	[15:0]	simplePinWrite_u423;
wire	[15:0]	simplePinWrite_u424;
wire		simplePinWrite_u425;
wire	[7:0]	simplePinWrite_u426;
wire	[15:0]	simplePinWrite_u427;
wire	[7:0]	simplePinWrite_u428;
wire		simplePinWrite_u429;
reg	[31:0]	syncEnable_u151=32'h0;
reg		reg_01db5434_u0=1'h0;
reg	[31:0]	syncEnable_u152_u0=32'h0;
reg		reg_014e92e3_u0=1'h0;
reg	[31:0]	syncEnable_u153_u0=32'h0;
assign add={port_01245fcb_[24:0], 7'b0}+{port_01245fcb_[26:0], 5'b0};
assign add_u561={add[31:5], 5'b0}+{port_01245fcb_[27:0], 4'b0};
assign add_u562={add_u561[31:4], 4'b0}+port_00c7b822_;
assign add_u563=32'h0+add_u562;
assign or_u363_u0=and_u1469_u0|RESET;
assign and_u1469_u0=done_cache_u16&port_012755fe_;
always @(posedge CLK or posedge reg_014e92e3_u0 or posedge or_u363_u0)
begin
if (or_u363_u0)
done_cache_u16<=1'h0;
else if (reg_014e92e3_u0)
done_cache_u16<=1'h1;
else done_cache_u16<=done_cache_u16;
end
assign add_u564={port_01245fcb_[24:0], 7'b0}+{port_01245fcb_[26:0], 5'b0};
assign add_u565={add_u564[31:5], 5'b0}+{port_01245fcb_[27:0], 4'b0};
assign add_u566={add_u565[31:4], 4'b0}+port_00c7b822_;
assign add_u567=32'h0+add_u566;
assign or_u364_u0=and_u1470_u0|RESET;
assign and_u1470_u0=done_cache_u17_u0&port_010e3311_;
always @(posedge CLK or posedge reg_014e92e3_u0 or posedge or_u364_u0)
begin
if (or_u364_u0)
done_cache_u17_u0<=1'h0;
else if (reg_014e92e3_u0)
done_cache_u17_u0<=1'h1;
else done_cache_u17_u0<=done_cache_u17_u0;
end
assign add_u568={port_01245fcb_[24:0], 7'b0}+{port_01245fcb_[26:0], 5'b0};
assign add_u569={add_u568[31:5], 5'b0}+{port_01245fcb_[27:0], 4'b0};
assign add_u570={add_u569[31:4], 4'b0}+port_00c7b822_;
assign add_u571=32'h0+add_u570;
assign and_u1471_u0=done_cache_u18_u0&port_00817c5e_;
assign or_u365_u0=and_u1471_u0|RESET;
always @(posedge CLK or posedge reg_014e92e3_u0 or posedge or_u365_u0)
begin
if (or_u365_u0)
done_cache_u18_u0<=1'h0;
else if (reg_014e92e3_u0)
done_cache_u18_u0<=1'h1;
else done_cache_u18_u0<=done_cache_u18_u0;
end
assign add_u572=port_00c7b822_+32'h1;
assign equals_a_signed=add_u572;
assign equals_b_signed=32'hb0;
assign equals=equals_a_signed==equals_b_signed;
assign and_u1472_u0=GO&not_u323_u0;
assign and_u1473_u0=GO&equals;
assign not_u323_u0=~equals;
assign add_u573=port_01245fcb_+32'h1;
assign mux_u262=(and_u1474_u0)?add_u572:32'h0;
assign and_u1474_u0=and_u1472_u0&GO;
assign and_u1475_u0=and_u1473_u0&GO;
assign mux_u263_u0=(and_u1474_u0)?port_01245fcb_:add_u573;
assign simplePinWrite=reg_01db5434_u0&{1{reg_01db5434_u0}};
assign simplePinWrite_u422=port_0041b215_;
assign simplePinWrite_u423=16'h1&{16{1'h1}};
assign simplePinWrite_u424=16'h1&{16{1'h1}};
assign simplePinWrite_u425=reg_01db5434_u0&{1{reg_01db5434_u0}};
assign simplePinWrite_u426=port_0148441b_;
assign simplePinWrite_u427=16'h1&{16{1'h1}};
assign simplePinWrite_u428=port_015914f6_;
assign simplePinWrite_u429=reg_01db5434_u0&{1{reg_01db5434_u0}};
always @(posedge CLK)
begin
if (GO)
syncEnable_u151<=add_u563;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01db5434_u0<=1'h0;
else reg_01db5434_u0<=reg_014e92e3_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u152_u0<=add_u571;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_014e92e3_u0<=1'h0;
else reg_014e92e3_u0<=GO;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u153_u0<=add_u567;
end
assign RESULT=GO;
assign RESULT_u1007=mux_u263_u0;
assign RESULT_u1008=GO;
assign RESULT_u1009=mux_u262;
assign RESULT_u1010=reg_014e92e3_u0;
assign RESULT_u1011=syncEnable_u152_u0;
assign RESULT_u1012=3'h1;
assign RESULT_u1013=reg_014e92e3_u0;
assign RESULT_u1014=syncEnable_u153_u0;
assign RESULT_u1015=3'h1;
assign RESULT_u1016=reg_014e92e3_u0;
assign RESULT_u1017=syncEnable_u151;
assign RESULT_u1018=3'h1;
assign RESULT_u1019=simplePinWrite_u422;
assign RESULT_u1020=simplePinWrite_u423;
assign RESULT_u1021=simplePinWrite_u424;
assign RESULT_u1022=simplePinWrite_u428;
assign RESULT_u1023=simplePinWrite;
assign RESULT_u1024=simplePinWrite_u429;
assign RESULT_u1025=simplePinWrite_u425;
assign RESULT_u1026=simplePinWrite_u427;
assign RESULT_u1027=simplePinWrite_u426;
assign DONE=reg_01db5434_u0;
endmodule



module PROCESS_stateVar_state_s1(bus_0008ca2f_, bus_0111fdbc_, bus_00e044d2_, bus_01b1cd40_, bus_0001e8b0_);
input		bus_0008ca2f_;
input		bus_0111fdbc_;
input		bus_00e044d2_;
input		bus_01b1cd40_;
output		bus_0001e8b0_;
reg		stateVar_state_s1_u19=1'h0;
always @(posedge bus_0008ca2f_ or posedge bus_0111fdbc_)
begin
if (bus_0111fdbc_)
stateVar_state_s1_u19<=1'h0;
else if (bus_00e044d2_)
stateVar_state_s1_u19<=bus_01b1cd40_;
end
assign bus_0001e8b0_=stateVar_state_s1_u19;
endmodule



module PROCESS_globalreset_physical_016c3655_(bus_00046cea_, bus_010f4e6e_, bus_01726b76_);
input		bus_00046cea_;
input		bus_010f4e6e_;
output		bus_01726b76_;
reg		sample_u34=1'h0;
reg		glitch_u34=1'h0;
wire		and_015cbb5e_u0;
reg		cross_u34=1'h0;
reg		final_u34=1'h1;
wire		or_01e64c9e_u0;
wire		not_00d23009_u0;
always @(posedge bus_00046cea_)
begin
sample_u34<=1'h1;
end
always @(posedge bus_00046cea_)
begin
glitch_u34<=cross_u34;
end
assign and_015cbb5e_u0=cross_u34&glitch_u34;
always @(posedge bus_00046cea_)
begin
cross_u34<=sample_u34;
end
always @(posedge bus_00046cea_)
begin
final_u34<=not_00d23009_u0;
end
assign bus_01726b76_=or_01e64c9e_u0;
assign or_01e64c9e_u0=bus_010f4e6e_|final_u34;
assign not_00d23009_u0=~and_015cbb5e_u0;
endmodule



module PROCESS_getValueRGB(CLK, RESET, GO, port_00285e4f_, port_00028fcf_, port_00612b21_, port_00100350_, port_01f41dbb_, port_0011132f_, port_00b6c0b7_, port_003f6d63_, RESULT, RESULT_u1028, RESULT_u1029, RESULT_u1030, RESULT_u1031, RESULT_u1032, RESULT_u1033, RESULT_u1034, RESULT_u1035, RESULT_u1036, RESULT_u1037, RESULT_u1038, RESULT_u1039, RESULT_u1040, RESULT_u1041, RESULT_u1042, RESULT_u1043, RESULT_u1044, RESULT_u1045, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_00285e4f_;
input	[31:0]	port_00028fcf_;
input		port_00612b21_;
input		port_00100350_;
input		port_01f41dbb_;
input	[7:0]	port_0011132f_;
input	[7:0]	port_00b6c0b7_;
input	[7:0]	port_003f6d63_;
output		RESULT;
output	[31:0]	RESULT_u1028;
output		RESULT_u1029;
output	[31:0]	RESULT_u1030;
output		RESULT_u1031;
output	[31:0]	RESULT_u1032;
output	[7:0]	RESULT_u1033;
output	[2:0]	RESULT_u1034;
output		RESULT_u1035;
output	[31:0]	RESULT_u1036;
output	[7:0]	RESULT_u1037;
output	[2:0]	RESULT_u1038;
output		RESULT_u1039;
output	[31:0]	RESULT_u1040;
output	[7:0]	RESULT_u1041;
output	[2:0]	RESULT_u1042;
output		RESULT_u1043;
output		RESULT_u1044;
output		RESULT_u1045;
output		DONE;
wire		simplePinWrite;
wire		simplePinWrite_u430;
wire		simplePinWrite_u431;
wire	[31:0]	add;
wire	[31:0]	add_u574;
wire	[31:0]	add_u575;
wire	[31:0]	add_u576;
wire		and_u1476_u0;
reg		reg_01694e95_u0=1'h0;
wire		or_u366_u0;
wire	[31:0]	add_u577;
wire	[31:0]	add_u578;
wire	[31:0]	add_u579;
wire	[31:0]	add_u580;
wire		and_u1477_u0;
wire		or_u367_u0;
reg		reg_01fde3c3_u0=1'h0;
wire	[31:0]	add_u581;
wire	[31:0]	add_u582;
wire	[31:0]	add_u583;
wire	[31:0]	add_u584;
reg		reg_01b9df05_u0=1'h0;
wire		or_u368_u0;
wire		and_u1478_u0;
wire	[31:0]	add_u585;
wire signed	[31:0]	equals_b_signed;
wire signed	[31:0]	equals_a_signed;
wire		equals;
wire		and_u1479_u0;
wire		and_u1480_u0;
wire		not_u324_u0;
wire	[31:0]	add_u586;
wire	[31:0]	mux_u264;
wire		and_u1481_u0;
wire		and_u1482_u0;
wire	[31:0]	mux_u265_u0;
reg	[7:0]	syncEnable_u154=8'h0;
reg	[7:0]	syncEnable_u155_u0=8'h0;
reg	[31:0]	syncEnable_u156_u0=32'h0;
reg		reg_01010ca3_u0=1'h0;
reg	[31:0]	syncEnable_u157_u0=32'h0;
reg	[7:0]	syncEnable_u158_u0=8'h0;
reg	[31:0]	syncEnable_u159_u0=32'h0;
reg		reg_01df0d3b_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign simplePinWrite_u430=GO&{1{GO}};
assign simplePinWrite_u431=GO&{1{GO}};
assign add={port_00285e4f_[24:0], 7'b0}+{port_00285e4f_[26:0], 5'b0};
assign add_u574={add[31:5], 5'b0}+{port_00285e4f_[27:0], 4'b0};
assign add_u575={add_u574[31:4], 4'b0}+port_00028fcf_;
assign add_u576=32'h0+add_u575;
assign and_u1476_u0=reg_01694e95_u0&port_01f41dbb_;
always @(posedge CLK or posedge reg_01df0d3b_u0 or posedge or_u366_u0)
begin
if (or_u366_u0)
reg_01694e95_u0<=1'h0;
else if (reg_01df0d3b_u0)
reg_01694e95_u0<=1'h1;
else reg_01694e95_u0<=reg_01694e95_u0;
end
assign or_u366_u0=and_u1476_u0|RESET;
assign add_u577={port_00285e4f_[24:0], 7'b0}+{port_00285e4f_[26:0], 5'b0};
assign add_u578={add_u577[31:5], 5'b0}+{port_00285e4f_[27:0], 4'b0};
assign add_u579={add_u578[31:4], 4'b0}+port_00028fcf_;
assign add_u580=32'h0+add_u579;
assign and_u1477_u0=reg_01fde3c3_u0&port_00100350_;
assign or_u367_u0=and_u1477_u0|RESET;
always @(posedge CLK or posedge reg_01df0d3b_u0 or posedge or_u367_u0)
begin
if (or_u367_u0)
reg_01fde3c3_u0<=1'h0;
else if (reg_01df0d3b_u0)
reg_01fde3c3_u0<=1'h1;
else reg_01fde3c3_u0<=reg_01fde3c3_u0;
end
assign add_u581={port_00285e4f_[24:0], 7'b0}+{port_00285e4f_[26:0], 5'b0};
assign add_u582={add_u581[31:5], 5'b0}+{port_00285e4f_[27:0], 4'b0};
assign add_u583={add_u582[31:4], 4'b0}+port_00028fcf_;
assign add_u584=32'h0+add_u583;
always @(posedge CLK or posedge reg_01df0d3b_u0 or posedge or_u368_u0)
begin
if (or_u368_u0)
reg_01b9df05_u0<=1'h0;
else if (reg_01df0d3b_u0)
reg_01b9df05_u0<=1'h1;
else reg_01b9df05_u0<=reg_01b9df05_u0;
end
assign or_u368_u0=and_u1478_u0|RESET;
assign and_u1478_u0=reg_01b9df05_u0&port_00612b21_;
assign add_u585=port_00028fcf_+32'h1;
assign equals_a_signed=add_u585;
assign equals_b_signed=32'hb0;
assign equals=equals_a_signed==equals_b_signed;
assign and_u1479_u0=GO&not_u324_u0;
assign and_u1480_u0=GO&equals;
assign not_u324_u0=~equals;
assign add_u586=port_00285e4f_+32'h1;
assign mux_u264=(and_u1482_u0)?32'h0:add_u585;
assign and_u1481_u0=and_u1479_u0&GO;
assign and_u1482_u0=and_u1480_u0&GO;
assign mux_u265_u0=(and_u1482_u0)?add_u586:port_00285e4f_;
always @(posedge CLK)
begin
if (GO)
syncEnable_u154<=port_003f6d63_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u155_u0<=port_00b6c0b7_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u156_u0<=add_u584;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01010ca3_u0<=1'h0;
else reg_01010ca3_u0<=reg_01df0d3b_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u157_u0<=add_u580;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u158_u0<=port_0011132f_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u159_u0<=add_u576;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01df0d3b_u0<=1'h0;
else reg_01df0d3b_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u1028=mux_u265_u0;
assign RESULT_u1029=GO;
assign RESULT_u1030=mux_u264;
assign RESULT_u1031=reg_01df0d3b_u0;
assign RESULT_u1032=syncEnable_u156_u0;
assign RESULT_u1033=syncEnable_u158_u0;
assign RESULT_u1034=3'h1;
assign RESULT_u1035=reg_01df0d3b_u0;
assign RESULT_u1036=syncEnable_u157_u0;
assign RESULT_u1037=syncEnable_u154;
assign RESULT_u1038=3'h1;
assign RESULT_u1039=reg_01df0d3b_u0;
assign RESULT_u1040=syncEnable_u159_u0;
assign RESULT_u1041=syncEnable_u155_u0;
assign RESULT_u1042=3'h1;
assign RESULT_u1043=simplePinWrite_u430;
assign RESULT_u1044=simplePinWrite_u431;
assign RESULT_u1045=simplePinWrite;
assign DONE=reg_01010ca3_u0;
endmodule



module PROCESS_simplememoryreferee_018cecb6_(bus_004bdde8_, bus_00d5e4f7_, bus_0074cb0b_, bus_0092b9ff_, bus_01655295_, bus_00ba52c3_, bus_0092895d_, bus_0018d135_, bus_00f11bd2_, bus_01a2f21a_, bus_010a585d_, bus_01a2e3de_, bus_017fc3a3_, bus_014f17a8_);
input		bus_004bdde8_;
input		bus_00d5e4f7_;
input		bus_0074cb0b_;
input	[7:0]	bus_0092b9ff_;
input		bus_01655295_;
input	[7:0]	bus_00ba52c3_;
input	[31:0]	bus_0092895d_;
input	[2:0]	bus_0018d135_;
output	[7:0]	bus_00f11bd2_;
output	[31:0]	bus_01a2f21a_;
output		bus_010a585d_;
output		bus_01a2e3de_;
output	[2:0]	bus_017fc3a3_;
output		bus_014f17a8_;
assign bus_00f11bd2_=8'hff;
assign bus_01a2f21a_=bus_0092895d_;
assign bus_010a585d_=bus_01655295_;
assign bus_01a2e3de_=bus_01655295_;
assign bus_017fc3a3_=3'h1;
assign bus_014f17a8_=bus_0074cb0b_;
endmodule



module PROCESS_simplememoryreferee_01df3566_(bus_00f883fe_, bus_01a1d096_, bus_01662e30_, bus_018b8df6_, bus_006e6d0c_, bus_00cc16ec_, bus_00dda92a_, bus_00381fab_, bus_01154382_, bus_013b413c_, bus_0166f79c_, bus_00e30286_, bus_015b67b7_, bus_00a7282d_);
input		bus_00f883fe_;
input		bus_01a1d096_;
input		bus_01662e30_;
input	[7:0]	bus_018b8df6_;
input		bus_006e6d0c_;
input	[7:0]	bus_00cc16ec_;
input	[31:0]	bus_00dda92a_;
input	[2:0]	bus_00381fab_;
output	[7:0]	bus_01154382_;
output	[31:0]	bus_013b413c_;
output		bus_0166f79c_;
output		bus_00e30286_;
output	[2:0]	bus_015b67b7_;
output		bus_00a7282d_;
assign bus_01154382_=8'h0;
assign bus_013b413c_=bus_00dda92a_;
assign bus_0166f79c_=bus_006e6d0c_;
assign bus_00e30286_=bus_006e6d0c_;
assign bus_015b67b7_=3'h1;
assign bus_00a7282d_=bus_01662e30_;
endmodule



module PROCESS_Kicker_34(CLK, RESET, bus_00709018_);
input		CLK;
input		RESET;
output		bus_00709018_;
wire		bus_013c8232_;
reg		kicker_1=1'h0;
reg		kicker_res=1'h0;
wire		bus_01d82959_;
reg		kicker_2=1'h0;
wire		bus_007cf3ae_;
wire		bus_014264db_;
assign bus_013c8232_=~RESET;
always @(posedge CLK)
begin
kicker_1<=bus_013c8232_;
end
always @(posedge CLK)
begin
kicker_res<=bus_01d82959_;
end
assign bus_01d82959_=kicker_1&bus_013c8232_&bus_007cf3ae_;
always @(posedge CLK)
begin
kicker_2<=bus_014264db_;
end
assign bus_007cf3ae_=~kicker_2;
assign bus_00709018_=kicker_res;
assign bus_014264db_=bus_013c8232_&kicker_1;
endmodule



module PROCESS_stateVar_state_s0(bus_01ae46ae_, bus_00a25ac8_, bus_000bdb25_, bus_0045f0e9_, bus_013a80a2_);
input		bus_01ae46ae_;
input		bus_00a25ac8_;
input		bus_000bdb25_;
input		bus_0045f0e9_;
output		bus_013a80a2_;
reg		stateVar_state_s0_u19=1'h0;
assign bus_013a80a2_=stateVar_state_s0_u19;
always @(posedge bus_01ae46ae_ or posedge bus_00a25ac8_)
begin
if (bus_00a25ac8_)
stateVar_state_s0_u19<=1'h0;
else if (bus_000bdb25_)
stateVar_state_s0_u19<=bus_0045f0e9_;
end
endmodule



module PROCESS_stateVar_state_s2(bus_01855671_, bus_00ee2f23_, bus_01cf20d2_, bus_01948536_, bus_0088e767_);
input		bus_01855671_;
input		bus_00ee2f23_;
input		bus_01cf20d2_;
input		bus_01948536_;
output		bus_0088e767_;
reg		stateVar_state_s2_u17=1'h0;
assign bus_0088e767_=stateVar_state_s2_u17;
always @(posedge bus_01855671_ or posedge bus_00ee2f23_)
begin
if (bus_00ee2f23_)
stateVar_state_s2_u17<=1'h0;
else if (bus_01cf20d2_)
stateVar_state_s2_u17<=bus_01948536_;
end
endmodule



module PROCESS_endianswapper_00f6c3f9_(endianswapper_00f6c3f9_in, endianswapper_00f6c3f9_out);
input	[31:0]	endianswapper_00f6c3f9_in;
output	[31:0]	endianswapper_00f6c3f9_out;
assign endianswapper_00f6c3f9_out=endianswapper_00f6c3f9_in;
endmodule



module PROCESS_endianswapper_019c5644_(endianswapper_019c5644_in, endianswapper_019c5644_out);
input	[31:0]	endianswapper_019c5644_in;
output	[31:0]	endianswapper_019c5644_out;
assign endianswapper_019c5644_out=endianswapper_019c5644_in;
endmodule



module PROCESS_stateVar_count_y(bus_01722449_, bus_00ac4f02_, bus_01303bc0_, bus_01483acc_, bus_0047b12a_, bus_01c6542c_, bus_009f3313_);
input		bus_01722449_;
input		bus_00ac4f02_;
input		bus_01303bc0_;
input	[31:0]	bus_01483acc_;
input		bus_0047b12a_;
input	[31:0]	bus_01c6542c_;
output	[31:0]	bus_009f3313_;
wire		or_0117e04e_u0;
reg	[31:0]	stateVar_count_y_u4=32'h0;
wire	[31:0]	mux_015a4e9c_u0;
wire	[31:0]	endianswapper_00f6c3f9_out;
wire	[31:0]	endianswapper_019c5644_out;
assign or_0117e04e_u0=bus_01303bc0_|bus_0047b12a_;
assign bus_009f3313_=endianswapper_00f6c3f9_out;
always @(posedge bus_01722449_ or posedge bus_00ac4f02_)
begin
if (bus_00ac4f02_)
stateVar_count_y_u4<=32'h0;
else if (or_0117e04e_u0)
stateVar_count_y_u4<=endianswapper_019c5644_out;
end
assign mux_015a4e9c_u0=(bus_01303bc0_)?bus_01483acc_:bus_01c6542c_;
PROCESS_endianswapper_00f6c3f9_ PROCESS_endianswapper_00f6c3f9__1(.endianswapper_00f6c3f9_in(stateVar_count_y_u4), 
  .endianswapper_00f6c3f9_out(endianswapper_00f6c3f9_out));
PROCESS_endianswapper_019c5644_ PROCESS_endianswapper_019c5644__1(.endianswapper_019c5644_in(mux_015a4e9c_u0), 
  .endianswapper_019c5644_out(endianswapper_019c5644_out));
endmodule



module PROCESS_simplememoryreferee_01e963df_(bus_00eb96d7_, bus_00fc372b_, bus_0123c590_, bus_00395682_, bus_007262df_, bus_00577cfe_, bus_004fde95_, bus_01289d14_, bus_005e8c9d_, bus_00a07c46_, bus_01ba61a9_, bus_0174247e_, bus_001f0d05_, bus_0160b5ac_);
input		bus_00eb96d7_;
input		bus_00fc372b_;
input		bus_0123c590_;
input	[7:0]	bus_00395682_;
input		bus_007262df_;
input	[7:0]	bus_00577cfe_;
input	[31:0]	bus_004fde95_;
input	[2:0]	bus_01289d14_;
output	[7:0]	bus_005e8c9d_;
output	[31:0]	bus_00a07c46_;
output		bus_01ba61a9_;
output		bus_0174247e_;
output	[2:0]	bus_001f0d05_;
output		bus_0160b5ac_;
assign bus_005e8c9d_=8'h0;
assign bus_00a07c46_=bus_004fde95_;
assign bus_01ba61a9_=bus_007262df_;
assign bus_0174247e_=bus_007262df_;
assign bus_001f0d05_=3'h1;
assign bus_0160b5ac_=bus_0123c590_;
endmodule



module PROCESS_structuralmemory_0145fced_(CLK_u18, bus_00ecf8c6_, bus_00703654_, bus_002a587c_, bus_012a3f30_, bus_00a4b4e9_, bus_01e65d20_, bus_00dfcb52_, bus_00d32323_, bus_00681dd1_, bus_006d22dd_, bus_009a9712_, bus_00ebe0d9_, bus_010bfe43_);
input		CLK_u18;
input		bus_00ecf8c6_;
input	[31:0]	bus_00703654_;
input	[2:0]	bus_002a587c_;
input		bus_012a3f30_;
input		bus_00a4b4e9_;
input	[7:0]	bus_01e65d20_;
input	[31:0]	bus_00dfcb52_;
input	[2:0]	bus_00d32323_;
input		bus_00681dd1_;
input	[7:0]	bus_006d22dd_;
output	[7:0]	bus_009a9712_;
output		bus_00ebe0d9_;
output		bus_010bfe43_;
reg		logicalMem_536c15_we_delay0_u0=1'h0;
wire	[7:0]	bus_00f9a8af_;
wire		or_01d2c323_u0;
reg		logicalMem_536c15_we_delay0_u1_u0=1'h0;
reg		logicalMem_536c15_re_delay0_u0=1'h0;
wire		or_019408d3_u0;
always @(posedge CLK_u18 or posedge bus_00ecf8c6_)
begin
if (bus_00ecf8c6_)
logicalMem_536c15_we_delay0_u0<=1'h0;
else logicalMem_536c15_we_delay0_u0<=bus_00a4b4e9_;
end
PROCESS_forge_memory_25344x8_27 PROCESS_forge_memory_25344x8_27_instance2(.CLK(CLK_u18), 
  .ENA(or_019408d3_u0), .WEA(bus_00a4b4e9_), .DINA(bus_01e65d20_), .ADDRA(bus_00703654_), 
  .DOUTA(bus_00f9a8af_), .DONEA(), .ENB(bus_00681dd1_), .WEB(bus_00681dd1_), .DINB(8'hff), 
  .ADDRB(bus_00dfcb52_), .DONEB());
assign or_01d2c323_u0=logicalMem_536c15_re_delay0_u0|logicalMem_536c15_we_delay0_u0;
assign bus_009a9712_=bus_00f9a8af_;
assign bus_00ebe0d9_=or_01d2c323_u0;
assign bus_010bfe43_=logicalMem_536c15_we_delay0_u1_u0;
always @(posedge CLK_u18 or posedge bus_00ecf8c6_)
begin
if (bus_00ecf8c6_)
logicalMem_536c15_we_delay0_u1_u0<=1'h0;
else logicalMem_536c15_we_delay0_u1_u0<=bus_00681dd1_;
end
always @(posedge CLK_u18 or posedge bus_00ecf8c6_)
begin
if (bus_00ecf8c6_)
logicalMem_536c15_re_delay0_u0<=1'h0;
else logicalMem_536c15_re_delay0_u0<=bus_012a3f30_;
end
assign or_019408d3_u0=bus_012a3f30_|bus_00a4b4e9_;
endmodule


