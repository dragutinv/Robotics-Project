// __  ___ __ ___  _ __   ___  ___ 
// \ \/ / '__/ _ \| '_ \ / _ \/ __|
//  >  <| | | (_) | | | | (_) \__ \
// /_/\_\_|  \___/|_| |_|\___/|___/
// 
// Xronos synthesizer version
// Run date: Wed 14 Oct 2015 15:56:36 +0100
// 

module output_process_Draw_rectangle(center_x_SEND, Gout_SEND, Bout_COUNT, Bin_SEND, Gin_SEND, center_y_ACK, Gout_RDY, Rin_COUNT, Rout_COUNT, Bout_RDY, center_y_COUNT, Gin_DATA, Gout_DATA, Bin_ACK, center_y_DATA, center_y_SEND, Bin_DATA, CLK, center_x_DATA, RESET, Bout_ACK, Gin_COUNT, Rout_RDY, center_x_ACK, center_x_COUNT, Rin_ACK, Gout_COUNT, Rin_SEND, Rout_DATA, Bout_DATA, Bin_COUNT, Bout_SEND, Rout_ACK, Gout_ACK, Rout_SEND, Gin_ACK, Rin_DATA);
wire		drawRectangle_go;
input		center_x_SEND;
wire		getCenterXY_go;
output		Gout_SEND;
wire		doneCountIm_go;
output	[15:0]	Bout_COUNT;
input		Bin_SEND;
input		Gin_SEND;
output		center_y_ACK;
input		Gout_RDY;
input	[15:0]	Rin_COUNT;
output	[15:0]	Rout_COUNT;
input		Bout_RDY;
wire		getValueRGB_done;
wire		doneCountIm_done;
input	[15:0]	center_y_COUNT;
input	[7:0]	Gin_DATA;
output	[7:0]	Gout_DATA;
output		Bin_ACK;
input	[15:0]	center_y_DATA;
input		center_y_SEND;
input	[7:0]	Bin_DATA;
input		CLK;
wire		getCenterXY_done;
input	[15:0]	center_x_DATA;
input		RESET;
input		Bout_ACK;
input	[15:0]	Gin_COUNT;
wire		send_done;
input		Rout_RDY;
output		center_x_ACK;
input	[15:0]	center_x_COUNT;
output		Rin_ACK;
output	[15:0]	Gout_COUNT;
wire		send_go;
input		Rin_SEND;
output	[7:0]	Rout_DATA;
output	[7:0]	Bout_DATA;
input	[15:0]	Bin_COUNT;
output		Bout_SEND;
input		Rout_ACK;
input		Gout_ACK;
output		Rout_SEND;
wire		getValueRGB_go;
wire		drawRectangle_done;
output		Gin_ACK;
input	[7:0]	Rin_DATA;
wire	[15:0]	bus_01d1a412_;
wire		bus_01077fcf_;
wire		bus_012c5118_;
wire	[7:0]	bus_00dfc9b7_;
wire	[31:0]	bus_00c286b0_;
wire	[2:0]	bus_011cb380_;
wire	[7:0]	bus_00d9fe67_;
wire		bus_0017baf9_;
wire		bus_01fdbc03_;
wire	[31:0]	bus_000450ed_;
wire		bus_006fd605_;
wire		bus_01c75ab7_;
wire		bus_010c1d9f_;
wire	[31:0]	bus_01b58b6c_;
wire		bus_00dca91e_;
wire		bus_00ce7b1d_;
wire	[31:0]	bus_00dd8deb_;
wire		bus_0111ea1a_;
wire		bus_00abd173_;
wire	[7:0]	bus_00b0eb42_;
wire	[7:0]	bus_00b899d0_;
wire		bus_001563a0_;
wire	[2:0]	bus_0179d231_;
wire		bus_00dadf33_;
wire		bus_0175ba82_;
wire		bus_0186ea08_;
wire	[2:0]	bus_002ee5f8_;
wire	[31:0]	bus_01c7605e_;
wire		bus_00cf6bd8_;
wire		bus_00a74b9d_;
wire	[7:0]	bus_00c8ef26_;
wire		bus_00f0fb51_;
wire		bus_005a91b0_;
wire	[7:0]	bus_0191448d_;
wire		output_process_Draw_rectangle_doneCountIm_instance_DONE;
wire		doneCountIm;
wire	[31:0]	doneCountIm_u7;
wire		bus_000768aa_;
wire	[2:0]	bus_00d2523f_;
wire	[7:0]	bus_00dfdcdb_;
wire		bus_004d7ac9_;
wire		bus_00222056_;
wire	[31:0]	bus_006317eb_;
wire		bus_00051f40_;
wire	[7:0]	bus_01bd6be1_;
wire		bus_01acb2ba_;
wire		bus_007bfbe5_;
wire	[7:0]	bus_01c4af42_;
wire		bus_01895947_;
wire		output_process_Draw_rectangle_send_instance_DONE;
wire	[31:0]	send_u110;
wire		send_u112;
wire		send_u109;
wire	[31:0]	send_u102;
wire	[7:0]	send_u115;
wire		send_u106;
wire	[7:0]	send_u114;
wire	[2:0]	send_u108;
wire	[15:0]	send_u120;
wire		send_u117;
wire		send_u103;
wire	[7:0]	send_u119;
wire	[15:0]	send_u118;
wire		send_u101;
wire	[2:0]	send_u111;
wire	[31:0]	send_u100;
wire	[31:0]	send_u104;
wire	[31:0]	send_u107;
wire		send;
wire	[15:0]	send_u116;
wire		send_u113;
wire	[2:0]	send_u105;
wire		bus_00826511_;
wire	[7:0]	drawRectangle_u28;
wire	[31:0]	drawRectangle_u43;
wire	[7:0]	drawRectangle_u36;
wire	[31:0]	drawRectangle_u39;
wire	[2:0]	drawRectangle_u29;
wire		drawRectangle_u34;
wire		drawRectangle_u42;
wire		drawRectangle_u38;
wire	[7:0]	drawRectangle_u44;
wire	[2:0]	drawRectangle_u33;
wire	[31:0]	drawRectangle_u31;
wire		drawRectangle_u30;
wire	[2:0]	drawRectangle_u25;
wire	[2:0]	drawRectangle_u41;
wire		output_process_Draw_rectangle_drawRectangle_instance_DONE;
wire	[31:0]	drawRectangle_u27;
wire	[31:0]	drawRectangle_u23;
wire	[31:0]	drawRectangle_u35;
wire	[2:0]	drawRectangle_u45;
wire	[7:0]	drawRectangle_u40;
wire	[7:0]	drawRectangle_u32;
wire	[7:0]	drawRectangle_u24;
wire	[2:0]	drawRectangle_u37;
wire		drawRectangle_u26;
wire		drawRectangle;
wire		getValueRGB;
wire	[31:0]	getValueRGB_u54;
wire	[7:0]	getValueRGB_u63;
wire		getValueRGB_u65;
wire	[31:0]	getValueRGB_u62;
wire		getValueRGB_u55;
wire		output_process_Draw_rectangle_getValueRGB_instance_DONE;
wire		getValueRGB_u70;
wire	[31:0]	getValueRGB_u66;
wire	[31:0]	getValueRGB_u56;
wire		getValueRGB_u71;
wire		getValueRGB_u57;
wire	[7:0]	getValueRGB_u59;
wire	[2:0]	getValueRGB_u60;
wire		getValueRGB_u61;
wire	[7:0]	getValueRGB_u67;
wire	[31:0]	getValueRGB_u58;
wire	[2:0]	getValueRGB_u64;
wire	[2:0]	getValueRGB_u68;
wire		getValueRGB_u69;
wire		bus_00e9d5a0_;
wire		bus_012a48ec_;
wire		bus_00c3bb80_;
wire		bus_01203b9e_;
wire	[7:0]	bus_008abdc8_;
wire		bus_00e4d935_;
wire	[31:0]	bus_015653dd_;
wire	[2:0]	bus_014758cb_;
wire		bus_015914b1_;
wire	[7:0]	bus_017f3e79_;
wire		bus_0119517f_;
wire	[15:0]	bus_01915a27_;
wire		bus_00eb1f11_;
wire		bus_0074d452_;
wire		bus_01ff134d_;
wire	[31:0]	bus_00b4f835_;
wire	[7:0]	bus_00a8f1e0_;
wire	[2:0]	bus_0076b457_;
wire		bus_008cf4be_;
wire		bus_0176022b_;
wire		bus_01cd028e_;
wire		scheduler_u239;
wire		scheduler;
wire		scheduler_u235;
wire		scheduler_u232;
wire		scheduler_u240;
wire		output_process_Draw_rectangle_scheduler_instance_DONE;
wire		scheduler_u241;
wire		scheduler_u238;
wire		scheduler_u231;
wire		scheduler_u237;
wire		scheduler_u234;
wire		scheduler_u233;
wire		scheduler_u230;
wire		scheduler_u236;
wire		bus_008215bb_;
wire		getCenterXY_u9;
wire		getCenterXY_u6;
wire	[15:0]	getCenterXY_u5;
wire		output_process_Draw_rectangle_getCenterXY_instance_DONE;
wire		getCenterXY;
wire		getCenterXY_u8;
wire	[15:0]	getCenterXY_u7;
assign drawRectangle_go=scheduler_u237;
assign getCenterXY_go=scheduler_u239;
assign Gout_SEND=send_u113;
assign doneCountIm_go=scheduler_u241;
assign Bout_COUNT=send_u116;
assign center_y_ACK=getCenterXY_u9;
assign Rout_COUNT=send_u118;
assign getValueRGB_done=bus_00eb1f11_;
assign doneCountIm_done=bus_01c75ab7_;
assign Gout_DATA=send_u119;
assign Bin_ACK=getValueRGB_u69;
assign getCenterXY_done=bus_012a48ec_;
assign send_done=bus_00dadf33_;
assign center_x_ACK=getCenterXY_u8;
assign Rin_ACK=getValueRGB_u71;
assign Gout_COUNT=send_u120;
assign send_go=scheduler_u238;
assign Rout_DATA=send_u114;
assign Bout_DATA=send_u115;
assign Bout_SEND=send_u117;
assign Rout_SEND=send_u112;
assign getValueRGB_go=scheduler_u240;
assign drawRectangle_done=bus_008215bb_;
assign Gin_ACK=getValueRGB_u70;
output_process_Draw_rectangle_stateVar_centre_x output_process_Draw_rectangle_stateVar_centre_x_1(.bus_00d7e567_(CLK), 
  .bus_0015fedc_(bus_00826511_), .bus_00f08bcd_(getCenterXY), .bus_00ee6ea9_(getCenterXY_u5), 
  .bus_01d1a412_(bus_01d1a412_));
output_process_Draw_rectangle_structuralmemory_0088abf5_ output_process_Draw_rectangle_structuralmemory_0088abf5__1(.CLK_u40(CLK), 
  .bus_01261a43_(bus_00826511_), .bus_012f92e5_(bus_01c7605e_), .bus_01a6b386_(3'h1), 
  .bus_0092d120_(bus_0186ea08_), .bus_00d0e113_(bus_00cf6bd8_), .bus_01ef33b7_(bus_0191448d_), 
  .bus_01fcf661_(bus_015653dd_), .bus_00f05729_(3'h1), .bus_01b7b159_(bus_00c3bb80_), 
  .bus_0085991d_(8'h0), .bus_00dfc9b7_(bus_00dfc9b7_), .bus_012c5118_(bus_012c5118_), 
  .bus_01077fcf_(bus_01077fcf_));
output_process_Draw_rectangle_stateVar_count_x output_process_Draw_rectangle_stateVar_count_x_1(.bus_006b286d_(CLK), 
  .bus_012b48d7_(bus_00826511_), .bus_0163cbd3_(getValueRGB), .bus_00445e9f_(getValueRGB_u54), 
  .bus_0089bc33_(doneCountIm), .bus_005f91d8_(32'h0), .bus_0168a5c8_(send), .bus_01719e1a_(send_u100), 
  .bus_00c286b0_(bus_00c286b0_));
output_process_Draw_rectangle_simplememoryreferee_00bd791e_ output_process_Draw_rectangle_simplememoryreferee_00bd791e__1(.bus_00f6e05a_(CLK), 
  .bus_00035501_(bus_00826511_), .bus_0000bc38_(bus_0119517f_), .bus_01ac44d1_(8'h0), 
  .bus_00bdd017_(drawRectangle_u38), .bus_01bbf55e_(8'hff), .bus_01497e84_(drawRectangle_u39), 
  .bus_01c87704_(3'h1), .bus_00d9fe67_(bus_00d9fe67_), .bus_000450ed_(bus_000450ed_), 
  .bus_0017baf9_(bus_0017baf9_), .bus_006fd605_(bus_006fd605_), .bus_011cb380_(bus_011cb380_), 
  .bus_01fdbc03_(bus_01fdbc03_));
assign bus_01c75ab7_=output_process_Draw_rectangle_doneCountIm_instance_DONE&{1{output_process_Draw_rectangle_doneCountIm_instance_DONE}};
output_process_Draw_rectangle_stateVar_state_s3 output_process_Draw_rectangle_stateVar_state_s3_1(.bus_0150cf6f_(CLK), 
  .bus_006296a0_(bus_00826511_), .bus_01f22cb1_(scheduler_u235), .bus_00a4709a_(scheduler_u236), 
  .bus_010c1d9f_(bus_010c1d9f_));
output_process_Draw_rectangle_stateVar_count_y output_process_Draw_rectangle_stateVar_count_y_1(.bus_0093d58b_(CLK), 
  .bus_01a8c307_(bus_00826511_), .bus_018bc5d9_(getValueRGB_u55), .bus_00526a03_(getValueRGB_u56), 
  .bus_00c8cb38_(send_u101), .bus_01ee9eff_(send_u102), .bus_01b58b6c_(bus_01b58b6c_));
output_process_Draw_rectangle_simplememoryreferee_00ed4e4b_ output_process_Draw_rectangle_simplememoryreferee_00ed4e4b__1(.bus_00986971_(CLK), 
  .bus_00329dec_(bus_00826511_), .bus_0176ddd4_(bus_015914b1_), .bus_00e281d0_(bus_017f3e79_), 
  .bus_01d9f95a_(getValueRGB_u61), .bus_009797a4_(getValueRGB_u63), .bus_00490a3d_(getValueRGB_u62), 
  .bus_0128a7a1_(3'h1), .bus_01aa6f62_(drawRectangle_u42), .bus_019d31a8_(8'hff), 
  .bus_00fcf048_(drawRectangle_u43), .bus_01fa2a04_(3'h1), .bus_01f34ea7_(send_u106), 
  .bus_015b02f8_(send_u107), .bus_01bc72c1_(3'h1), .bus_00b899d0_(bus_00b899d0_), 
  .bus_00dd8deb_(bus_00dd8deb_), .bus_00ce7b1d_(bus_00ce7b1d_), .bus_00abd173_(bus_00abd173_), 
  .bus_0179d231_(bus_0179d231_), .bus_001563a0_(bus_001563a0_), .bus_00dca91e_(bus_00dca91e_), 
  .bus_00b0eb42_(bus_00b0eb42_), .bus_0111ea1a_(bus_0111ea1a_));
assign bus_00dadf33_=output_process_Draw_rectangle_send_instance_DONE&{1{output_process_Draw_rectangle_send_instance_DONE}};
output_process_Draw_rectangle_stateVar_state_s1 output_process_Draw_rectangle_stateVar_state_s1_1(.bus_0026e8e4_(CLK), 
  .bus_0083eb7b_(bus_00826511_), .bus_01d89dfc_(scheduler_u231), .bus_01aa2d2b_(scheduler_u232), 
  .bus_0175ba82_(bus_0175ba82_));
output_process_Draw_rectangle_simplememoryreferee_00e73508_ output_process_Draw_rectangle_simplememoryreferee_00e73508__1(.bus_0097f1ee_(CLK), 
  .bus_018c70c6_(bus_00826511_), .bus_005ad139_(bus_012c5118_), .bus_0097d2cf_(bus_00dfc9b7_), 
  .bus_01379b18_(getValueRGB_u65), .bus_01f860ed_(getValueRGB_u67), .bus_014410c3_(getValueRGB_u66), 
  .bus_0119f9bb_(3'h1), .bus_000c8909_(drawRectangle), .bus_00d8cc3c_(8'h0), .bus_00513dc1_(drawRectangle_u23), 
  .bus_00cb5bb1_(3'h1), .bus_018a06de_(send_u103), .bus_01e5a8d9_(send_u104), .bus_006aefd4_(3'h1), 
  .bus_0191448d_(bus_0191448d_), .bus_01c7605e_(bus_01c7605e_), .bus_00cf6bd8_(bus_00cf6bd8_), 
  .bus_0186ea08_(bus_0186ea08_), .bus_002ee5f8_(bus_002ee5f8_), .bus_005a91b0_(bus_005a91b0_), 
  .bus_00f0fb51_(bus_00f0fb51_), .bus_00c8ef26_(bus_00c8ef26_), .bus_00a74b9d_(bus_00a74b9d_));
output_process_Draw_rectangle_doneCountIm output_process_Draw_rectangle_doneCountIm_instance(.CLK(CLK), 
  .RESET(bus_00826511_), .GO(doneCountIm_go), .RESULT(doneCountIm), .RESULT_u1005(doneCountIm_u7), 
  .DONE(output_process_Draw_rectangle_doneCountIm_instance_DONE));
output_process_Draw_rectangle_simplememoryreferee_00b19833_ output_process_Draw_rectangle_simplememoryreferee_00b19833__1(.bus_014864e4_(CLK), 
  .bus_01d7d21d_(bus_00826511_), .bus_01cdbc0b_(bus_01895947_), .bus_00731aba_(bus_01c4af42_), 
  .bus_00c05064_(getValueRGB_u57), .bus_016bbcb6_(getValueRGB_u59), .bus_00d1ab4d_(getValueRGB_u58), 
  .bus_014bf606_(3'h1), .bus_00ae72f1_(drawRectangle_u26), .bus_00a8c929_(8'h0), 
  .bus_0090b74f_(drawRectangle_u27), .bus_015a01a5_(3'h1), .bus_00e606a1_(send_u109), 
  .bus_01d3e50a_(send_u110), .bus_00f86e25_(3'h1), .bus_00dfdcdb_(bus_00dfdcdb_), 
  .bus_006317eb_(bus_006317eb_), .bus_01acb2ba_(bus_01acb2ba_), .bus_004d7ac9_(bus_004d7ac9_), 
  .bus_00d2523f_(bus_00d2523f_), .bus_00051f40_(bus_00051f40_), .bus_00222056_(bus_00222056_), 
  .bus_01bd6be1_(bus_01bd6be1_), .bus_000768aa_(bus_000768aa_));
output_process_Draw_rectangle_structuralmemory_009e6b31_ output_process_Draw_rectangle_structuralmemory_009e6b31__1(.CLK_u41(CLK), 
  .bus_00b032dc_(bus_00826511_), .bus_01964486_(bus_006317eb_), .bus_0028847c_(3'h1), 
  .bus_01184a86_(bus_004d7ac9_), .bus_00d02e4c_(bus_01acb2ba_), .bus_00a2e19a_(bus_00dfdcdb_), 
  .bus_0024fc7c_(bus_00b4f835_), .bus_011d5d2a_(3'h1), .bus_006c78c2_(bus_01ff134d_), 
  .bus_012c686d_(8'h0), .bus_01c4af42_(bus_01c4af42_), .bus_01895947_(bus_01895947_), 
  .bus_007bfbe5_(bus_007bfbe5_));
output_process_Draw_rectangle_send output_process_Draw_rectangle_send_instance(.CLK(CLK), 
  .RESET(bus_00826511_), .GO(send_go), .port_0002ea05_(bus_00c286b0_), .port_002f724a_(bus_01b58b6c_), 
  .port_0125acd4_(bus_00a74b9d_), .port_002687bf_(bus_00c8ef26_), .port_000fa29b_(bus_0111ea1a_), 
  .port_00f9e1da_(bus_00b0eb42_), .port_0038b572_(bus_000768aa_), .port_0122d684_(bus_01bd6be1_), 
  .RESULT(send), .RESULT_u1006(send_u100), .RESULT_u1007(send_u101), .RESULT_u1008(send_u102), 
  .RESULT_u1015(send_u103), .RESULT_u1016(send_u104), .RESULT_u1017(send_u105), 
  .RESULT_u1009(send_u106), .RESULT_u1010(send_u107), .RESULT_u1011(send_u108), 
  .RESULT_u1012(send_u109), .RESULT_u1013(send_u110), .RESULT_u1014(send_u111), 
  .RESULT_u1018(send_u112), .RESULT_u1019(send_u113), .RESULT_u1021(send_u114), 
  .RESULT_u1020(send_u115), .RESULT_u1022(send_u116), .RESULT_u1023(send_u117), 
  .RESULT_u1024(send_u118), .RESULT_u1026(send_u119), .RESULT_u1025(send_u120), 
  .DONE(output_process_Draw_rectangle_send_instance_DONE));
output_process_Draw_rectangle_globalreset_physical_001fa2b7_ output_process_Draw_rectangle_globalreset_physical_001fa2b7__1(.bus_0023db22_(CLK), 
  .bus_0113813a_(RESET), .bus_00826511_(bus_00826511_));
output_process_Draw_rectangle_drawRectangle output_process_Draw_rectangle_drawRectangle_instance(.CLK(CLK), 
  .RESET(bus_00826511_), .GO(drawRectangle_go), .port_00be099f_(bus_01915a27_), 
  .port_0116e071_(bus_01d1a412_), .port_01a2503a_(bus_00f0fb51_), .port_01d67dc6_(bus_00222056_), 
  .port_018e9e2f_(bus_0176022b_), .port_0087f92c_(bus_01203b9e_), .port_00891739_(bus_01fdbc03_), 
  .port_000bb648_(bus_00dca91e_), .RESULT_u1034(drawRectangle), .RESULT_u1035(drawRectangle_u23), 
  .RESULT_u1036(drawRectangle_u24), .RESULT_u1037(drawRectangle_u25), .RESULT_u1030(drawRectangle_u26), 
  .RESULT_u1031(drawRectangle_u27), .RESULT_u1032(drawRectangle_u28), .RESULT_u1033(drawRectangle_u29), 
  .RESULT_u1046(drawRectangle_u30), .RESULT_u1047(drawRectangle_u31), .RESULT_u1048(drawRectangle_u32), 
  .RESULT_u1049(drawRectangle_u33), .RESULT_u1042(drawRectangle_u34), .RESULT_u1043(drawRectangle_u35), 
  .RESULT_u1044(drawRectangle_u36), .RESULT_u1045(drawRectangle_u37), .RESULT_u1038(drawRectangle_u38), 
  .RESULT_u1039(drawRectangle_u39), .RESULT_u1040(drawRectangle_u40), .RESULT_u1041(drawRectangle_u41), 
  .RESULT(drawRectangle_u42), .RESULT_u1027(drawRectangle_u43), .RESULT_u1028(drawRectangle_u44), 
  .RESULT_u1029(drawRectangle_u45), .DONE(output_process_Draw_rectangle_drawRectangle_instance_DONE));
output_process_Draw_rectangle_getValueRGB output_process_Draw_rectangle_getValueRGB_instance(.CLK(CLK), 
  .RESET(bus_00826511_), .GO(getValueRGB_go), .port_00c91e9e_(bus_00c286b0_), .port_00c1d6b4_(bus_01b58b6c_), 
  .port_01e0f363_(bus_00051f40_), .port_00aa595c_(bus_001563a0_), .port_006e1316_(bus_005a91b0_), 
  .port_016b104e_(Bin_DATA), .port_00a96b61_(Rin_DATA), .port_004f15e5_(Gin_DATA), 
  .RESULT(getValueRGB), .RESULT_u1050(getValueRGB_u54), .RESULT_u1051(getValueRGB_u55), 
  .RESULT_u1052(getValueRGB_u56), .RESULT_u1057(getValueRGB_u57), .RESULT_u1058(getValueRGB_u58), 
  .RESULT_u1059(getValueRGB_u59), .RESULT_u1060(getValueRGB_u60), .RESULT_u1053(getValueRGB_u61), 
  .RESULT_u1054(getValueRGB_u62), .RESULT_u1055(getValueRGB_u63), .RESULT_u1056(getValueRGB_u64), 
  .RESULT_u1061(getValueRGB_u65), .RESULT_u1062(getValueRGB_u66), .RESULT_u1063(getValueRGB_u67), 
  .RESULT_u1064(getValueRGB_u68), .RESULT_u1065(getValueRGB_u69), .RESULT_u1066(getValueRGB_u70), 
  .RESULT_u1067(getValueRGB_u71), .DONE(output_process_Draw_rectangle_getValueRGB_instance_DONE));
output_process_Draw_rectangle_Kicker_21 output_process_Draw_rectangle_Kicker_21_1(.CLK(CLK), 
  .RESET(bus_00826511_), .bus_00e9d5a0_(bus_00e9d5a0_));
assign bus_012a48ec_=output_process_Draw_rectangle_getCenterXY_instance_DONE&{1{output_process_Draw_rectangle_getCenterXY_instance_DONE}};
output_process_Draw_rectangle_simplememoryreferee_01bc888a_ output_process_Draw_rectangle_simplememoryreferee_01bc888a__1(.bus_00150c03_(CLK), 
  .bus_01c7b9d3_(bus_00826511_), .bus_01179579_(bus_01077fcf_), .bus_01764864_(8'h0), 
  .bus_00a40f07_(drawRectangle_u34), .bus_00bb1f5c_(8'h0), .bus_010d3878_(drawRectangle_u35), 
  .bus_002943c5_(3'h1), .bus_008abdc8_(bus_008abdc8_), .bus_015653dd_(bus_015653dd_), 
  .bus_00c3bb80_(bus_00c3bb80_), .bus_00e4d935_(bus_00e4d935_), .bus_014758cb_(bus_014758cb_), 
  .bus_01203b9e_(bus_01203b9e_));
output_process_Draw_rectangle_structuralmemory_0198cbd9_ output_process_Draw_rectangle_structuralmemory_0198cbd9__1(.CLK_u42(CLK), 
  .bus_01d301f6_(bus_00826511_), .bus_01c3d072_(bus_00dd8deb_), .bus_014da5cc_(3'h1), 
  .bus_0169c6de_(bus_00abd173_), .bus_014ecd16_(bus_00ce7b1d_), .bus_01437b60_(bus_00b899d0_), 
  .bus_01e5c110_(bus_000450ed_), .bus_00c30c8e_(3'h1), .bus_0143d8b1_(bus_0017baf9_), 
  .bus_0031ac17_(8'hff), .bus_017f3e79_(bus_017f3e79_), .bus_015914b1_(bus_015914b1_), 
  .bus_0119517f_(bus_0119517f_));
output_process_Draw_rectangle_stateVar_centre_y output_process_Draw_rectangle_stateVar_centre_y_1(.bus_008068bf_(CLK), 
  .bus_005cd3da_(bus_00826511_), .bus_002324b9_(getCenterXY_u6), .bus_00e92383_(getCenterXY_u7), 
  .bus_01915a27_(bus_01915a27_));
assign bus_00eb1f11_=output_process_Draw_rectangle_getValueRGB_instance_DONE&{1{output_process_Draw_rectangle_getValueRGB_instance_DONE}};
output_process_Draw_rectangle_stateVar_state_s0 output_process_Draw_rectangle_stateVar_state_s0_1(.bus_012cd072_(CLK), 
  .bus_01290bbe_(bus_00826511_), .bus_00c0ada5_(scheduler), .bus_002ce97c_(scheduler_u230), 
  .bus_0074d452_(bus_0074d452_));
output_process_Draw_rectangle_simplememoryreferee_00d7a4d7_ output_process_Draw_rectangle_simplememoryreferee_00d7a4d7__1(.bus_0121612e_(CLK), 
  .bus_00732c35_(bus_00826511_), .bus_009da5d7_(bus_007bfbe5_), .bus_005076d2_(8'h0), 
  .bus_0188d17c_(drawRectangle_u30), .bus_0138f3bb_(8'h0), .bus_01d679a0_(drawRectangle_u31), 
  .bus_00aa30fc_(3'h1), .bus_00a8f1e0_(bus_00a8f1e0_), .bus_00b4f835_(bus_00b4f835_), 
  .bus_01ff134d_(bus_01ff134d_), .bus_008cf4be_(bus_008cf4be_), .bus_0076b457_(bus_0076b457_), 
  .bus_0176022b_(bus_0176022b_));
output_process_Draw_rectangle_stateVar_state_s2 output_process_Draw_rectangle_stateVar_state_s2_1(.bus_00f238fa_(CLK), 
  .bus_007ac458_(bus_00826511_), .bus_005d6340_(scheduler_u233), .bus_000dff53_(scheduler_u234), 
  .bus_01cd028e_(bus_01cd028e_));
output_process_Draw_rectangle_scheduler output_process_Draw_rectangle_scheduler_instance(.CLK(CLK), 
  .RESET(bus_00826511_), .GO(bus_00e9d5a0_), .port_003e9bda_(bus_0074d452_), .port_01961eea_(bus_0175ba82_), 
  .port_0012bfe7_(bus_01cd028e_), .port_0055998f_(bus_010c1d9f_), .port_01f67390_(bus_00c286b0_), 
  .port_000bbff8_(center_x_SEND), .port_01b61592_(getCenterXY_done), .port_0091ced8_(doneCountIm_done), 
  .port_002e8e34_(Rin_SEND), .port_01613518_(Bin_SEND), .port_0192ec25_(Gin_SEND), 
  .port_01ca5227_(center_y_SEND), .port_01559388_(Rout_RDY), .port_00cb09f8_(send_done), 
  .port_01572c5f_(Gout_RDY), .port_012d89fe_(drawRectangle_done), .port_009db78a_(Bout_RDY), 
  .port_007e9851_(getValueRGB_done), .RESULT(scheduler), .RESULT_u1068(scheduler_u230), 
  .RESULT_u1069(scheduler_u231), .RESULT_u1070(scheduler_u232), .RESULT_u1071(scheduler_u233), 
  .RESULT_u1072(scheduler_u234), .RESULT_u1073(scheduler_u235), .RESULT_u1074(scheduler_u236), 
  .RESULT_u1076(scheduler_u237), .RESULT_u1075(scheduler_u238), .RESULT_u1077(scheduler_u239), 
  .RESULT_u1079(scheduler_u240), .RESULT_u1078(scheduler_u241), .DONE(output_process_Draw_rectangle_scheduler_instance_DONE));
assign bus_008215bb_=output_process_Draw_rectangle_drawRectangle_instance_DONE&{1{output_process_Draw_rectangle_drawRectangle_instance_DONE}};
output_process_Draw_rectangle_getCenterXY output_process_Draw_rectangle_getCenterXY_instance(.CLK(CLK), 
  .RESET(bus_00826511_), .GO(getCenterXY_go), .port_002f348e_(center_y_DATA), .port_0163315b_(center_x_DATA), 
  .RESULT(getCenterXY), .RESULT_u1080(getCenterXY_u5), .RESULT_u1081(getCenterXY_u6), 
  .RESULT_u1082(getCenterXY_u7), .RESULT_u1083(getCenterXY_u8), .RESULT_u1084(getCenterXY_u9), 
  .DONE(output_process_Draw_rectangle_getCenterXY_instance_DONE));
endmodule



module output_process_Draw_rectangle_endianswapper_0089b0f2_(endianswapper_0089b0f2_in, endianswapper_0089b0f2_out);
input	[15:0]	endianswapper_0089b0f2_in;
output	[15:0]	endianswapper_0089b0f2_out;
assign endianswapper_0089b0f2_out=endianswapper_0089b0f2_in;
endmodule



module output_process_Draw_rectangle_endianswapper_00593a7d_(endianswapper_00593a7d_in, endianswapper_00593a7d_out);
input	[15:0]	endianswapper_00593a7d_in;
output	[15:0]	endianswapper_00593a7d_out;
assign endianswapper_00593a7d_out=endianswapper_00593a7d_in;
endmodule



module output_process_Draw_rectangle_stateVar_centre_x(bus_00d7e567_, bus_0015fedc_, bus_00f08bcd_, bus_00ee6ea9_, bus_01d1a412_);
input		bus_00d7e567_;
input		bus_0015fedc_;
input		bus_00f08bcd_;
input	[15:0]	bus_00ee6ea9_;
output	[15:0]	bus_01d1a412_;
reg	[15:0]	stateVar_centre_x_u5=16'h0;
wire	[15:0]	endianswapper_0089b0f2_out;
wire	[15:0]	endianswapper_00593a7d_out;
assign bus_01d1a412_=endianswapper_00593a7d_out;
always @(posedge bus_00d7e567_ or posedge bus_0015fedc_)
begin
if (bus_0015fedc_)
stateVar_centre_x_u5<=16'h0;
else if (bus_00f08bcd_)
stateVar_centre_x_u5<=endianswapper_0089b0f2_out;
end
output_process_Draw_rectangle_endianswapper_0089b0f2_ output_process_Draw_rectangle_endianswapper_0089b0f2__1(.endianswapper_0089b0f2_in(bus_00ee6ea9_), 
  .endianswapper_0089b0f2_out(endianswapper_0089b0f2_out));
output_process_Draw_rectangle_endianswapper_00593a7d_ output_process_Draw_rectangle_endianswapper_00593a7d__1(.endianswapper_00593a7d_in(stateVar_centre_x_u5), 
  .endianswapper_00593a7d_out(endianswapper_00593a7d_out));
endmodule



module output_process_Draw_rectangle_forge_memory_25344x8_69(CLK, ENA, WEA, DINA, ENB, WEB, DINB, ADDRA, ADDRB, DOUTA, DONEA, DONEB);
input		CLK;
input		ENA;
input		WEA;
input	[7:0]	DINA;
input		ENB;
input		WEB;
input	[7:0]	DINB;
input	[31:0]	ADDRA;
input	[31:0]	ADDRB;
output	[7:0]	DOUTA;
output		DONEA;
output		DONEB;
wire		wea_0;
wire		web_0;
wire	[7:0]	pre_douta_0;
wire		wea_1;
wire		web_1;
wire	[7:0]	pre_douta_1;
reg	[7:0]	mux_outa;
reg	[31:0]	ADDRA_reg;
reg	[31:0]	ADDRB_reg;
wire	[7:0]	pre_doutb_0;
reg	[7:0]	mux_outb;
wire	[7:0]	pre_doutb_1;
reg		web_done;
reg		rea_done;
reg		wea_done;
assign wea_0=WEA&(ADDRA[31:14]==18'h0);
assign web_0=WEB&(ADDRB[31:14]==18'h0);
assign wea_1=WEA&(ADDRA[31:14]==18'h1);
assign web_1=WEB&(ADDRB[31:14]==18'h1);
always @(posedge CLK)
begin
ADDRA_reg<=ADDRA;
end
always @(ADDRA_reg or pre_douta_0 or pre_douta_1)
begin
case (ADDRA_reg[31:14])18'd0:mux_outa=pre_douta_0;
18'd1:mux_outa=pre_douta_1;
default:mux_outa=8'h0;
endcase end
always @(posedge CLK)
begin
ADDRB_reg<=ADDRB;
end
always @(ADDRB_reg or pre_doutb_0 or pre_doutb_1)
begin
case (ADDRB_reg[31:14])18'd0:mux_outb=pre_doutb_0;
18'd1:mux_outb=pre_doutb_1;
default:mux_outb=8'h0;
endcase end
always @(posedge CLK)
begin
wea_done<=WEA;
rea_done<=ENA;
web_done<=WEB;
end
assign DONEA=wea_done|rea_done;
assign DONEB=web_done;
assign DOUTA=mux_outa;
// Memory array element: COL: 0, ROW: 0
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_72(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[0]), .DOA(pre_douta_0[0]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[0]), .DOB());
// Memory array element: COL: 0, ROW: 1
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_73(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[1]), .DOA(pre_douta_0[1]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[1]), .DOB());
// Memory array element: COL: 0, ROW: 2
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_74(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[2]), .DOA(pre_douta_0[2]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[2]), .DOB());
// Memory array element: COL: 0, ROW: 3
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_75(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[3]), .DOA(pre_douta_0[3]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[3]), .DOB());
// Memory array element: COL: 0, ROW: 4
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_76(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[4]), .DOA(pre_douta_0[4]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[4]), .DOB());
// Memory array element: COL: 0, ROW: 5
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_77(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[5]), .DOA(pre_douta_0[5]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[5]), .DOB());
// Memory array element: COL: 0, ROW: 6
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_78(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[6]), .DOA(pre_douta_0[6]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[6]), .DOB());
// Memory array element: COL: 0, ROW: 7
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_79(.CLKA(CLK), 
  .WEA(wea_0), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[7]), .DOA(pre_douta_0[7]), 
  .CLKB(CLK), .WEB(web_0), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[7]), .DOB());
// Memory array element: COL: 1, ROW: 0
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_80(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[0]), .DOA(pre_douta_1[0]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[0]), .DOB());
// Memory array element: COL: 1, ROW: 1
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_81(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[1]), .DOA(pre_douta_1[1]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[1]), .DOB());
// Memory array element: COL: 1, ROW: 2
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_82(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[2]), .DOA(pre_douta_1[2]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[2]), .DOB());
// Memory array element: COL: 1, ROW: 3
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_83(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[3]), .DOA(pre_douta_1[3]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[3]), .DOB());
// Memory array element: COL: 1, ROW: 4
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_84(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[4]), .DOA(pre_douta_1[4]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[4]), .DOB());
// Memory array element: COL: 1, ROW: 5
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_85(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[5]), .DOA(pre_douta_1[5]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[5]), .DOB());
// Memory array element: COL: 1, ROW: 6
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_86(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[6]), .DOA(pre_douta_1[6]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[6]), .DOB());
// Memory array element: COL: 1, ROW: 7
//  Initialization of Dual Port Block ram now done through explicit
// parameter setting.
RAMB16_S1_S1#(.INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000), 
  .WRITE_MODE_A("READ_FIRST"), .WRITE_MODE_B("READ_FIRST"))RAMB16_S1_S1_instance_87(.CLKA(CLK), 
  .WEA(wea_1), .ENA(ENA), .SSRA(1'b0), .ADDRA(ADDRA), .DIA(DINA[7]), .DOA(pre_douta_1[7]), 
  .CLKB(CLK), .WEB(web_1), .ENB(ENB), .SSRB(1'b0), .ADDRB(ADDRB), .DIB(DINB[7]), .DOB());
endmodule



module output_process_Draw_rectangle_structuralmemory_0088abf5_(CLK_u40, bus_01261a43_, bus_012f92e5_, bus_01a6b386_, bus_0092d120_, bus_00d0e113_, bus_01ef33b7_, bus_01fcf661_, bus_00f05729_, bus_01b7b159_, bus_0085991d_, bus_00dfc9b7_, bus_012c5118_, bus_01077fcf_);
input		CLK_u40;
input		bus_01261a43_;
input	[31:0]	bus_012f92e5_;
input	[2:0]	bus_01a6b386_;
input		bus_0092d120_;
input		bus_00d0e113_;
input	[7:0]	bus_01ef33b7_;
input	[31:0]	bus_01fcf661_;
input	[2:0]	bus_00f05729_;
input		bus_01b7b159_;
input	[7:0]	bus_0085991d_;
output	[7:0]	bus_00dfc9b7_;
output		bus_012c5118_;
output		bus_01077fcf_;
reg		logicalMem_c35a43_we_delay0_u0=1'h0;
reg		logicalMem_c35a43_we_delay0_u1_u0=1'h0;
wire		or_01592923_u0;
wire	[7:0]	bus_00ef53af_;
wire		or_010a4259_u0;
reg		logicalMem_c35a43_re_delay0_u0=1'h0;
always @(posedge CLK_u40 or posedge bus_01261a43_)
begin
if (bus_01261a43_)
logicalMem_c35a43_we_delay0_u0<=1'h0;
else logicalMem_c35a43_we_delay0_u0<=bus_01b7b159_;
end
always @(posedge CLK_u40 or posedge bus_01261a43_)
begin
if (bus_01261a43_)
logicalMem_c35a43_we_delay0_u1_u0<=1'h0;
else logicalMem_c35a43_we_delay0_u1_u0<=bus_00d0e113_;
end
assign or_01592923_u0=logicalMem_c35a43_re_delay0_u0|logicalMem_c35a43_we_delay0_u1_u0;
output_process_Draw_rectangle_forge_memory_25344x8_69 output_process_Draw_rectangle_forge_memory_25344x8_69_instance0(.CLK(CLK_u40), 
  .ENA(or_010a4259_u0), .WEA(bus_00d0e113_), .DINA(bus_01ef33b7_), .ADDRA(bus_012f92e5_), 
  .DOUTA(bus_00ef53af_), .DONEA(), .ENB(bus_01b7b159_), .WEB(bus_01b7b159_), .DINB(8'h0), 
  .ADDRB(bus_01fcf661_), .DONEB());
assign or_010a4259_u0=bus_0092d120_|bus_00d0e113_;
assign bus_00dfc9b7_=bus_00ef53af_;
assign bus_012c5118_=or_01592923_u0;
assign bus_01077fcf_=logicalMem_c35a43_we_delay0_u0;
always @(posedge CLK_u40 or posedge bus_01261a43_)
begin
if (bus_01261a43_)
logicalMem_c35a43_re_delay0_u0<=1'h0;
else logicalMem_c35a43_re_delay0_u0<=bus_0092d120_;
end
endmodule



module output_process_Draw_rectangle_endianswapper_00295635_(endianswapper_00295635_in, endianswapper_00295635_out);
input	[31:0]	endianswapper_00295635_in;
output	[31:0]	endianswapper_00295635_out;
assign endianswapper_00295635_out=endianswapper_00295635_in;
endmodule



module output_process_Draw_rectangle_endianswapper_002ab668_(endianswapper_002ab668_in, endianswapper_002ab668_out);
input	[31:0]	endianswapper_002ab668_in;
output	[31:0]	endianswapper_002ab668_out;
assign endianswapper_002ab668_out=endianswapper_002ab668_in;
endmodule



module output_process_Draw_rectangle_stateVar_count_x(bus_006b286d_, bus_012b48d7_, bus_0163cbd3_, bus_00445e9f_, bus_0089bc33_, bus_005f91d8_, bus_0168a5c8_, bus_01719e1a_, bus_00c286b0_);
input		bus_006b286d_;
input		bus_012b48d7_;
input		bus_0163cbd3_;
input	[31:0]	bus_00445e9f_;
input		bus_0089bc33_;
input	[31:0]	bus_005f91d8_;
input		bus_0168a5c8_;
input	[31:0]	bus_01719e1a_;
output	[31:0]	bus_00c286b0_;
wire	[31:0]	endianswapper_00295635_out;
wire	[31:0]	endianswapper_002ab668_out;
wire		or_019fa15c_u0;
wire	[31:0]	mux_01aed992_u0;
reg	[31:0]	stateVar_count_x_u7=32'h0;
output_process_Draw_rectangle_endianswapper_00295635_ output_process_Draw_rectangle_endianswapper_00295635__1(.endianswapper_00295635_in(mux_01aed992_u0), 
  .endianswapper_00295635_out(endianswapper_00295635_out));
output_process_Draw_rectangle_endianswapper_002ab668_ output_process_Draw_rectangle_endianswapper_002ab668__1(.endianswapper_002ab668_in(stateVar_count_x_u7), 
  .endianswapper_002ab668_out(endianswapper_002ab668_out));
assign or_019fa15c_u0=bus_0163cbd3_|bus_0089bc33_|bus_0168a5c8_;
assign mux_01aed992_u0=({32{bus_0163cbd3_}}&bus_00445e9f_)|({32{bus_0089bc33_}}&32'h0)|({32{bus_0168a5c8_}}&bus_01719e1a_);
always @(posedge bus_006b286d_ or posedge bus_012b48d7_)
begin
if (bus_012b48d7_)
stateVar_count_x_u7<=32'h0;
else if (or_019fa15c_u0)
stateVar_count_x_u7<=endianswapper_00295635_out;
end
assign bus_00c286b0_=endianswapper_002ab668_out;
endmodule



module output_process_Draw_rectangle_simplememoryreferee_00bd791e_(bus_00f6e05a_, bus_00035501_, bus_0000bc38_, bus_01ac44d1_, bus_00bdd017_, bus_01bbf55e_, bus_01497e84_, bus_01c87704_, bus_00d9fe67_, bus_000450ed_, bus_0017baf9_, bus_006fd605_, bus_011cb380_, bus_01fdbc03_);
input		bus_00f6e05a_;
input		bus_00035501_;
input		bus_0000bc38_;
input	[7:0]	bus_01ac44d1_;
input		bus_00bdd017_;
input	[7:0]	bus_01bbf55e_;
input	[31:0]	bus_01497e84_;
input	[2:0]	bus_01c87704_;
output	[7:0]	bus_00d9fe67_;
output	[31:0]	bus_000450ed_;
output		bus_0017baf9_;
output		bus_006fd605_;
output	[2:0]	bus_011cb380_;
output		bus_01fdbc03_;
assign bus_00d9fe67_=8'hff;
assign bus_000450ed_=bus_01497e84_;
assign bus_0017baf9_=bus_00bdd017_;
assign bus_006fd605_=bus_00bdd017_;
assign bus_011cb380_=3'h1;
assign bus_01fdbc03_=bus_0000bc38_;
endmodule



module output_process_Draw_rectangle_stateVar_state_s3(bus_0150cf6f_, bus_006296a0_, bus_01f22cb1_, bus_00a4709a_, bus_010c1d9f_);
input		bus_0150cf6f_;
input		bus_006296a0_;
input		bus_01f22cb1_;
input		bus_00a4709a_;
output		bus_010c1d9f_;
reg		stateVar_state_s3_u10=1'h0;
assign bus_010c1d9f_=stateVar_state_s3_u10;
always @(posedge bus_0150cf6f_ or posedge bus_006296a0_)
begin
if (bus_006296a0_)
stateVar_state_s3_u10<=1'h0;
else if (bus_01f22cb1_)
stateVar_state_s3_u10<=bus_00a4709a_;
end
endmodule



module output_process_Draw_rectangle_endianswapper_00e87db1_(endianswapper_00e87db1_in, endianswapper_00e87db1_out);
input	[31:0]	endianswapper_00e87db1_in;
output	[31:0]	endianswapper_00e87db1_out;
assign endianswapper_00e87db1_out=endianswapper_00e87db1_in;
endmodule



module output_process_Draw_rectangle_endianswapper_018c8696_(endianswapper_018c8696_in, endianswapper_018c8696_out);
input	[31:0]	endianswapper_018c8696_in;
output	[31:0]	endianswapper_018c8696_out;
assign endianswapper_018c8696_out=endianswapper_018c8696_in;
endmodule



module output_process_Draw_rectangle_stateVar_count_y(bus_0093d58b_, bus_01a8c307_, bus_018bc5d9_, bus_00526a03_, bus_00c8cb38_, bus_01ee9eff_, bus_01b58b6c_);
input		bus_0093d58b_;
input		bus_01a8c307_;
input		bus_018bc5d9_;
input	[31:0]	bus_00526a03_;
input		bus_00c8cb38_;
input	[31:0]	bus_01ee9eff_;
output	[31:0]	bus_01b58b6c_;
reg	[31:0]	stateVar_count_y_u7=32'h0;
wire	[31:0]	mux_00bb7e3a_u0;
wire		or_0125ffb1_u0;
wire	[31:0]	endianswapper_00e87db1_out;
wire	[31:0]	endianswapper_018c8696_out;
always @(posedge bus_0093d58b_ or posedge bus_01a8c307_)
begin
if (bus_01a8c307_)
stateVar_count_y_u7<=32'h0;
else if (or_0125ffb1_u0)
stateVar_count_y_u7<=endianswapper_018c8696_out;
end
assign mux_00bb7e3a_u0=(bus_018bc5d9_)?bus_00526a03_:bus_01ee9eff_;
assign or_0125ffb1_u0=bus_018bc5d9_|bus_00c8cb38_;
assign bus_01b58b6c_=endianswapper_00e87db1_out;
output_process_Draw_rectangle_endianswapper_00e87db1_ output_process_Draw_rectangle_endianswapper_00e87db1__1(.endianswapper_00e87db1_in(stateVar_count_y_u7), 
  .endianswapper_00e87db1_out(endianswapper_00e87db1_out));
output_process_Draw_rectangle_endianswapper_018c8696_ output_process_Draw_rectangle_endianswapper_018c8696__1(.endianswapper_018c8696_in(mux_00bb7e3a_u0), 
  .endianswapper_018c8696_out(endianswapper_018c8696_out));
endmodule



module output_process_Draw_rectangle_simplememoryreferee_00ed4e4b_(bus_00986971_, bus_00329dec_, bus_0176ddd4_, bus_00e281d0_, bus_01d9f95a_, bus_009797a4_, bus_00490a3d_, bus_0128a7a1_, bus_01aa6f62_, bus_019d31a8_, bus_00fcf048_, bus_01fa2a04_, bus_01f34ea7_, bus_015b02f8_, bus_01bc72c1_, bus_00b899d0_, bus_00dd8deb_, bus_00ce7b1d_, bus_00abd173_, bus_0179d231_, bus_001563a0_, bus_00dca91e_, bus_00b0eb42_, bus_0111ea1a_);
input		bus_00986971_;
input		bus_00329dec_;
input		bus_0176ddd4_;
input	[7:0]	bus_00e281d0_;
input		bus_01d9f95a_;
input	[7:0]	bus_009797a4_;
input	[31:0]	bus_00490a3d_;
input	[2:0]	bus_0128a7a1_;
input		bus_01aa6f62_;
input	[7:0]	bus_019d31a8_;
input	[31:0]	bus_00fcf048_;
input	[2:0]	bus_01fa2a04_;
input		bus_01f34ea7_;
input	[31:0]	bus_015b02f8_;
input	[2:0]	bus_01bc72c1_;
output	[7:0]	bus_00b899d0_;
output	[31:0]	bus_00dd8deb_;
output		bus_00ce7b1d_;
output		bus_00abd173_;
output	[2:0]	bus_0179d231_;
output		bus_001563a0_;
output		bus_00dca91e_;
output	[7:0]	bus_00b0eb42_;
output		bus_0111ea1a_;
wire		not_01e2a94c_u0;
wire		or_00d8302e_u0;
wire		or_01b8ea2c_u0;
reg		done_qual_u83=1'h0;
wire		or_00c4afbc_u0;
wire		or_00c68761_u0;
reg		done_qual_u84_u0=1'h0;
wire	[31:0]	mux_01e644e2_u0;
wire		and_019dfb4e_u0;
wire		and_0188eef3_u0;
wire		not_009b6a17_u0;
reg		done_qual_u85_u0=1'h0;
wire		not_00b7e754_u0;
wire		and_00ecd6c8_u0;
wire	[7:0]	mux_014035d6_u0;
wire		or_01c68acc_u0;
assign not_01e2a94c_u0=~bus_0176ddd4_;
assign or_00d8302e_u0=bus_01d9f95a_|bus_01aa6f62_;
assign or_01b8ea2c_u0=bus_01d9f95a_|done_qual_u85_u0;
always @(posedge bus_00986971_)
begin
if (bus_00329dec_)
done_qual_u83<=1'h0;
else done_qual_u83<=bus_01f34ea7_;
end
assign or_00c4afbc_u0=bus_01aa6f62_|done_qual_u84_u0;
assign or_00c68761_u0=bus_01f34ea7_|done_qual_u83;
always @(posedge bus_00986971_)
begin
if (bus_00329dec_)
done_qual_u84_u0<=1'h0;
else done_qual_u84_u0<=bus_01aa6f62_;
end
assign bus_00b899d0_=mux_014035d6_u0;
assign bus_00dd8deb_=mux_01e644e2_u0;
assign bus_00ce7b1d_=or_00d8302e_u0;
assign bus_00abd173_=or_01c68acc_u0;
assign bus_0179d231_=3'h1;
assign bus_001563a0_=and_00ecd6c8_u0;
assign bus_00dca91e_=and_0188eef3_u0;
assign bus_00b0eb42_=bus_00e281d0_;
assign bus_0111ea1a_=and_019dfb4e_u0;
assign mux_01e644e2_u0=({32{bus_01d9f95a_}}&bus_00490a3d_)|({32{bus_01aa6f62_}}&bus_00fcf048_)|({32{bus_01f34ea7_}}&bus_015b02f8_);
assign and_019dfb4e_u0=or_00c68761_u0&bus_0176ddd4_;
assign and_0188eef3_u0=or_00c4afbc_u0&bus_0176ddd4_;
assign not_009b6a17_u0=~bus_0176ddd4_;
always @(posedge bus_00986971_)
begin
if (bus_00329dec_)
done_qual_u85_u0<=1'h0;
else done_qual_u85_u0<=bus_01d9f95a_;
end
assign not_00b7e754_u0=~bus_0176ddd4_;
assign and_00ecd6c8_u0=or_01b8ea2c_u0&bus_0176ddd4_;
assign mux_014035d6_u0=(bus_01d9f95a_)?bus_009797a4_:8'hff;
assign or_01c68acc_u0=bus_01d9f95a_|bus_01aa6f62_|bus_01f34ea7_;
endmodule



module output_process_Draw_rectangle_stateVar_state_s1(bus_0026e8e4_, bus_0083eb7b_, bus_01d89dfc_, bus_01aa2d2b_, bus_0175ba82_);
input		bus_0026e8e4_;
input		bus_0083eb7b_;
input		bus_01d89dfc_;
input		bus_01aa2d2b_;
output		bus_0175ba82_;
reg		stateVar_state_s1_u18=1'h0;
assign bus_0175ba82_=stateVar_state_s1_u18;
always @(posedge bus_0026e8e4_ or posedge bus_0083eb7b_)
begin
if (bus_0083eb7b_)
stateVar_state_s1_u18<=1'h0;
else if (bus_01d89dfc_)
stateVar_state_s1_u18<=bus_01aa2d2b_;
end
endmodule



module output_process_Draw_rectangle_simplememoryreferee_00e73508_(bus_0097f1ee_, bus_018c70c6_, bus_005ad139_, bus_0097d2cf_, bus_01379b18_, bus_01f860ed_, bus_014410c3_, bus_0119f9bb_, bus_000c8909_, bus_00d8cc3c_, bus_00513dc1_, bus_00cb5bb1_, bus_018a06de_, bus_01e5a8d9_, bus_006aefd4_, bus_0191448d_, bus_01c7605e_, bus_00cf6bd8_, bus_0186ea08_, bus_002ee5f8_, bus_005a91b0_, bus_00f0fb51_, bus_00c8ef26_, bus_00a74b9d_);
input		bus_0097f1ee_;
input		bus_018c70c6_;
input		bus_005ad139_;
input	[7:0]	bus_0097d2cf_;
input		bus_01379b18_;
input	[7:0]	bus_01f860ed_;
input	[31:0]	bus_014410c3_;
input	[2:0]	bus_0119f9bb_;
input		bus_000c8909_;
input	[7:0]	bus_00d8cc3c_;
input	[31:0]	bus_00513dc1_;
input	[2:0]	bus_00cb5bb1_;
input		bus_018a06de_;
input	[31:0]	bus_01e5a8d9_;
input	[2:0]	bus_006aefd4_;
output	[7:0]	bus_0191448d_;
output	[31:0]	bus_01c7605e_;
output		bus_00cf6bd8_;
output		bus_0186ea08_;
output	[2:0]	bus_002ee5f8_;
output		bus_005a91b0_;
output		bus_00f0fb51_;
output	[7:0]	bus_00c8ef26_;
output		bus_00a74b9d_;
wire		or_01aa7fe1_u0;
wire		not_00a47ffe_u0;
wire		and_0113c05f_u0;
wire		and_0083fcff_u0;
wire		or_0049c916_u0;
wire		or_01b2f0d3_u0;
reg		done_qual_u86_u0=1'h0;
reg		done_qual_u87_u0=1'h0;
wire		or_014c9556_u0;
wire		not_01de481d_u0;
reg		done_qual_u88_u0=1'h0;
wire		or_01fafe59_u0;
wire	[31:0]	mux_000cc7c7_u0;
wire	[7:0]	mux_00b002d3_u0;
wire		and_0016924b_u0;
wire		not_0051fcaa_u0;
assign or_01aa7fe1_u0=bus_01379b18_|bus_000c8909_|bus_018a06de_;
assign not_00a47ffe_u0=~bus_005ad139_;
assign and_0113c05f_u0=or_0049c916_u0&bus_005ad139_;
assign and_0083fcff_u0=or_01b2f0d3_u0&bus_005ad139_;
assign or_0049c916_u0=bus_01379b18_|done_qual_u86_u0;
assign or_01b2f0d3_u0=bus_000c8909_|done_qual_u88_u0;
always @(posedge bus_0097f1ee_)
begin
if (bus_018c70c6_)
done_qual_u86_u0<=1'h0;
else done_qual_u86_u0<=bus_01379b18_;
end
always @(posedge bus_0097f1ee_)
begin
if (bus_018c70c6_)
done_qual_u87_u0<=1'h0;
else done_qual_u87_u0<=bus_018a06de_;
end
assign or_014c9556_u0=bus_01379b18_|bus_000c8909_;
assign not_01de481d_u0=~bus_005ad139_;
always @(posedge bus_0097f1ee_)
begin
if (bus_018c70c6_)
done_qual_u88_u0<=1'h0;
else done_qual_u88_u0<=bus_000c8909_;
end
assign or_01fafe59_u0=bus_018a06de_|done_qual_u87_u0;
assign mux_000cc7c7_u0=({32{bus_01379b18_}}&bus_014410c3_)|({32{bus_000c8909_}}&bus_00513dc1_)|({32{bus_018a06de_}}&bus_01e5a8d9_);
assign mux_00b002d3_u0=(bus_01379b18_)?bus_01f860ed_:8'h0;
assign and_0016924b_u0=or_01fafe59_u0&bus_005ad139_;
assign not_0051fcaa_u0=~bus_005ad139_;
assign bus_0191448d_=mux_00b002d3_u0;
assign bus_01c7605e_=mux_000cc7c7_u0;
assign bus_00cf6bd8_=or_014c9556_u0;
assign bus_0186ea08_=or_01aa7fe1_u0;
assign bus_002ee5f8_=3'h1;
assign bus_005a91b0_=and_0113c05f_u0;
assign bus_00f0fb51_=and_0083fcff_u0;
assign bus_00c8ef26_=bus_0097d2cf_;
assign bus_00a74b9d_=and_0016924b_u0;
endmodule



module output_process_Draw_rectangle_doneCountIm(CLK, RESET, GO, RESULT, RESULT_u1005, DONE);
input		CLK;
input		RESET;
input		GO;
output		RESULT;
output	[31:0]	RESULT_u1005;
output		DONE;
reg		reg_01549e55_u0=1'h0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01549e55_u0<=1'h0;
else reg_01549e55_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u1005=32'h0;
assign DONE=reg_01549e55_u0;
endmodule



module output_process_Draw_rectangle_simplememoryreferee_00b19833_(bus_014864e4_, bus_01d7d21d_, bus_01cdbc0b_, bus_00731aba_, bus_00c05064_, bus_016bbcb6_, bus_00d1ab4d_, bus_014bf606_, bus_00ae72f1_, bus_00a8c929_, bus_0090b74f_, bus_015a01a5_, bus_00e606a1_, bus_01d3e50a_, bus_00f86e25_, bus_00dfdcdb_, bus_006317eb_, bus_01acb2ba_, bus_004d7ac9_, bus_00d2523f_, bus_00051f40_, bus_00222056_, bus_01bd6be1_, bus_000768aa_);
input		bus_014864e4_;
input		bus_01d7d21d_;
input		bus_01cdbc0b_;
input	[7:0]	bus_00731aba_;
input		bus_00c05064_;
input	[7:0]	bus_016bbcb6_;
input	[31:0]	bus_00d1ab4d_;
input	[2:0]	bus_014bf606_;
input		bus_00ae72f1_;
input	[7:0]	bus_00a8c929_;
input	[31:0]	bus_0090b74f_;
input	[2:0]	bus_015a01a5_;
input		bus_00e606a1_;
input	[31:0]	bus_01d3e50a_;
input	[2:0]	bus_00f86e25_;
output	[7:0]	bus_00dfdcdb_;
output	[31:0]	bus_006317eb_;
output		bus_01acb2ba_;
output		bus_004d7ac9_;
output	[2:0]	bus_00d2523f_;
output		bus_00051f40_;
output		bus_00222056_;
output	[7:0]	bus_01bd6be1_;
output		bus_000768aa_;
wire		or_01f383d0_u0;
reg		done_qual_u89_u0=1'h0;
wire		or_00a848e4_u0;
wire		not_01804356_u0;
wire		or_0135612e_u0;
wire	[7:0]	mux_0037bc7d_u0;
reg		done_qual_u90_u0=1'h0;
wire		and_0072f1c6_u0;
wire		not_01027f4e_u0;
wire		or_0131a2c4_u0;
wire	[31:0]	mux_01c42324_u0;
reg		done_qual_u91_u0=1'h0;
wire		or_00ccd55d_u0;
wire		and_0033bbde_u0;
wire		not_00146daa_u0;
wire		and_019b4e25_u0;
assign or_01f383d0_u0=bus_00c05064_|bus_00ae72f1_;
always @(posedge bus_014864e4_)
begin
if (bus_01d7d21d_)
done_qual_u89_u0<=1'h0;
else done_qual_u89_u0<=bus_00c05064_;
end
assign bus_00dfdcdb_=mux_0037bc7d_u0;
assign bus_006317eb_=mux_01c42324_u0;
assign bus_01acb2ba_=or_01f383d0_u0;
assign bus_004d7ac9_=or_0131a2c4_u0;
assign bus_00d2523f_=3'h1;
assign bus_00051f40_=and_0033bbde_u0;
assign bus_00222056_=and_0072f1c6_u0;
assign bus_01bd6be1_=bus_00731aba_;
assign bus_000768aa_=and_019b4e25_u0;
assign or_00a848e4_u0=bus_00c05064_|done_qual_u89_u0;
assign not_01804356_u0=~bus_01cdbc0b_;
assign or_0135612e_u0=bus_00ae72f1_|done_qual_u91_u0;
assign mux_0037bc7d_u0=(bus_00c05064_)?bus_016bbcb6_:8'h0;
always @(posedge bus_014864e4_)
begin
if (bus_01d7d21d_)
done_qual_u90_u0<=1'h0;
else done_qual_u90_u0<=bus_00e606a1_;
end
assign and_0072f1c6_u0=or_0135612e_u0&bus_01cdbc0b_;
assign not_01027f4e_u0=~bus_01cdbc0b_;
assign or_0131a2c4_u0=bus_00c05064_|bus_00ae72f1_|bus_00e606a1_;
assign mux_01c42324_u0=({32{bus_00c05064_}}&bus_00d1ab4d_)|({32{bus_00ae72f1_}}&bus_0090b74f_)|({32{bus_00e606a1_}}&bus_01d3e50a_);
always @(posedge bus_014864e4_)
begin
if (bus_01d7d21d_)
done_qual_u91_u0<=1'h0;
else done_qual_u91_u0<=bus_00ae72f1_;
end
assign or_00ccd55d_u0=bus_00e606a1_|done_qual_u90_u0;
assign and_0033bbde_u0=or_00a848e4_u0&bus_01cdbc0b_;
assign not_00146daa_u0=~bus_01cdbc0b_;
assign and_019b4e25_u0=or_00ccd55d_u0&bus_01cdbc0b_;
endmodule



module output_process_Draw_rectangle_structuralmemory_009e6b31_(CLK_u41, bus_00b032dc_, bus_01964486_, bus_0028847c_, bus_01184a86_, bus_00d02e4c_, bus_00a2e19a_, bus_0024fc7c_, bus_011d5d2a_, bus_006c78c2_, bus_012c686d_, bus_01c4af42_, bus_01895947_, bus_007bfbe5_);
input		CLK_u41;
input		bus_00b032dc_;
input	[31:0]	bus_01964486_;
input	[2:0]	bus_0028847c_;
input		bus_01184a86_;
input		bus_00d02e4c_;
input	[7:0]	bus_00a2e19a_;
input	[31:0]	bus_0024fc7c_;
input	[2:0]	bus_011d5d2a_;
input		bus_006c78c2_;
input	[7:0]	bus_012c686d_;
output	[7:0]	bus_01c4af42_;
output		bus_01895947_;
output		bus_007bfbe5_;
wire		or_001822f1_u0;
reg		logicalMem_cc186b_re_delay0_u0=1'h0;
reg		logicalMem_cc186b_we_delay0_u0=1'h0;
reg		logicalMem_cc186b_we_delay0_u1_u0=1'h0;
wire		or_00f3bb30_u0;
wire	[7:0]	bus_016587e1_;
assign or_001822f1_u0=logicalMem_cc186b_re_delay0_u0|logicalMem_cc186b_we_delay0_u0;
always @(posedge CLK_u41 or posedge bus_00b032dc_)
begin
if (bus_00b032dc_)
logicalMem_cc186b_re_delay0_u0<=1'h0;
else logicalMem_cc186b_re_delay0_u0<=bus_01184a86_;
end
always @(posedge CLK_u41 or posedge bus_00b032dc_)
begin
if (bus_00b032dc_)
logicalMem_cc186b_we_delay0_u0<=1'h0;
else logicalMem_cc186b_we_delay0_u0<=bus_00d02e4c_;
end
always @(posedge CLK_u41 or posedge bus_00b032dc_)
begin
if (bus_00b032dc_)
logicalMem_cc186b_we_delay0_u1_u0<=1'h0;
else logicalMem_cc186b_we_delay0_u1_u0<=bus_006c78c2_;
end
assign bus_01c4af42_=bus_016587e1_;
assign bus_01895947_=or_001822f1_u0;
assign bus_007bfbe5_=logicalMem_cc186b_we_delay0_u1_u0;
assign or_00f3bb30_u0=bus_01184a86_|bus_00d02e4c_;
output_process_Draw_rectangle_forge_memory_25344x8_69 output_process_Draw_rectangle_forge_memory_25344x8_69_instance1(.CLK(CLK_u41), 
  .ENA(or_00f3bb30_u0), .WEA(bus_00d02e4c_), .DINA(bus_00a2e19a_), .ADDRA(bus_01964486_), 
  .DOUTA(bus_016587e1_), .DONEA(), .ENB(bus_006c78c2_), .WEB(bus_006c78c2_), .DINB(8'h0), 
  .ADDRB(bus_0024fc7c_), .DONEB());
endmodule



module output_process_Draw_rectangle_send(CLK, RESET, GO, port_0002ea05_, port_002f724a_, port_000fa29b_, port_00f9e1da_, port_0038b572_, port_0122d684_, port_0125acd4_, port_002687bf_, RESULT, RESULT_u1006, RESULT_u1007, RESULT_u1008, RESULT_u1009, RESULT_u1010, RESULT_u1011, RESULT_u1012, RESULT_u1013, RESULT_u1014, RESULT_u1015, RESULT_u1016, RESULT_u1017, RESULT_u1018, RESULT_u1019, RESULT_u1020, RESULT_u1021, RESULT_u1022, RESULT_u1023, RESULT_u1024, RESULT_u1025, RESULT_u1026, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_0002ea05_;
input	[31:0]	port_002f724a_;
input		port_000fa29b_;
input	[7:0]	port_00f9e1da_;
input		port_0038b572_;
input	[7:0]	port_0122d684_;
input		port_0125acd4_;
input	[7:0]	port_002687bf_;
output		RESULT;
output	[31:0]	RESULT_u1006;
output		RESULT_u1007;
output	[31:0]	RESULT_u1008;
output		RESULT_u1009;
output	[31:0]	RESULT_u1010;
output	[2:0]	RESULT_u1011;
output		RESULT_u1012;
output	[31:0]	RESULT_u1013;
output	[2:0]	RESULT_u1014;
output		RESULT_u1015;
output	[31:0]	RESULT_u1016;
output	[2:0]	RESULT_u1017;
output		RESULT_u1018;
output		RESULT_u1019;
output	[7:0]	RESULT_u1020;
output	[7:0]	RESULT_u1021;
output	[15:0]	RESULT_u1022;
output		RESULT_u1023;
output	[15:0]	RESULT_u1024;
output	[15:0]	RESULT_u1025;
output	[7:0]	RESULT_u1026;
output		DONE;
wire	[31:0]	add;
wire	[31:0]	add_u462;
wire	[31:0]	add_u463;
wire	[31:0]	add_u464;
wire		and_u1572_u0;
reg		done_cache_u54=1'h0;
wire		or_u434_u0;
wire	[31:0]	add_u465;
wire	[31:0]	add_u466;
wire	[31:0]	add_u467;
wire	[31:0]	add_u468;
wire		or_u435_u0;
wire		and_u1573_u0;
reg		done_cache_u55_u0=1'h0;
wire	[31:0]	add_u469;
wire	[31:0]	add_u470;
wire	[31:0]	add_u471;
wire	[31:0]	add_u472;
reg		done_cache_u56_u0=1'h0;
wire		and_u1574_u0;
wire		or_u436_u0;
wire	[31:0]	add_u473;
wire signed	[31:0]	equals_a_signed;
wire		equals;
wire signed	[31:0]	equals_b_signed;
wire		and_u1575_u0;
wire		and_u1576_u0;
wire		not_u325_u0;
wire	[31:0]	add_u474;
wire		and_u1577_u0;
wire		and_u1578_u0;
wire	[31:0]	mux_u498;
wire	[31:0]	mux_u499_u0;
wire		simplePinWrite;
wire	[7:0]	simplePinWrite_u237;
wire	[15:0]	simplePinWrite_u238;
wire	[15:0]	simplePinWrite_u239;
wire	[7:0]	simplePinWrite_u240;
wire		simplePinWrite_u241;
wire		simplePinWrite_u242;
wire	[15:0]	simplePinWrite_u243;
wire	[7:0]	simplePinWrite_u244;
reg	[31:0]	syncEnable_u360=32'h0;
reg	[31:0]	syncEnable_u361_u0=32'h0;
reg		reg_00b48d11_u0=1'h0;
reg		reg_013422da_u0=1'h0;
reg	[31:0]	syncEnable_u362_u0=32'h0;
assign add={port_0002ea05_[24:0], 7'b0}+{port_0002ea05_[26:0], 5'b0};
assign add_u462={add[31:5], 5'b0}+{port_0002ea05_[27:0], 4'b0};
assign add_u463={add_u462[31:4], 4'b0}+port_002f724a_;
assign add_u464=32'h0+add_u463;
assign and_u1572_u0=done_cache_u54&port_000fa29b_;
always @(posedge CLK or posedge reg_013422da_u0 or posedge or_u434_u0)
begin
if (or_u434_u0)
done_cache_u54<=1'h0;
else if (reg_013422da_u0)
done_cache_u54<=1'h1;
else done_cache_u54<=done_cache_u54;
end
assign or_u434_u0=and_u1572_u0|RESET;
assign add_u465={port_0002ea05_[24:0], 7'b0}+{port_0002ea05_[26:0], 5'b0};
assign add_u466={add_u465[31:5], 5'b0}+{port_0002ea05_[27:0], 4'b0};
assign add_u467={add_u466[31:4], 4'b0}+port_002f724a_;
assign add_u468=32'h0+add_u467;
assign or_u435_u0=and_u1573_u0|RESET;
assign and_u1573_u0=done_cache_u55_u0&port_0038b572_;
always @(posedge CLK or posedge reg_013422da_u0 or posedge or_u435_u0)
begin
if (or_u435_u0)
done_cache_u55_u0<=1'h0;
else if (reg_013422da_u0)
done_cache_u55_u0<=1'h1;
else done_cache_u55_u0<=done_cache_u55_u0;
end
assign add_u469={port_0002ea05_[24:0], 7'b0}+{port_0002ea05_[26:0], 5'b0};
assign add_u470={add_u469[31:5], 5'b0}+{port_0002ea05_[27:0], 4'b0};
assign add_u471={add_u470[31:4], 4'b0}+port_002f724a_;
assign add_u472=32'h0+add_u471;
always @(posedge CLK or posedge reg_013422da_u0 or posedge or_u436_u0)
begin
if (or_u436_u0)
done_cache_u56_u0<=1'h0;
else if (reg_013422da_u0)
done_cache_u56_u0<=1'h1;
else done_cache_u56_u0<=done_cache_u56_u0;
end
assign and_u1574_u0=done_cache_u56_u0&port_0125acd4_;
assign or_u436_u0=and_u1574_u0|RESET;
assign add_u473=port_002f724a_+32'h1;
assign equals_a_signed=add_u473;
assign equals_b_signed=32'hb0;
assign equals=equals_a_signed==equals_b_signed;
assign and_u1575_u0=GO&equals;
assign and_u1576_u0=GO&not_u325_u0;
assign not_u325_u0=~equals;
assign add_u474=port_0002ea05_+32'h1;
assign and_u1577_u0=and_u1575_u0&GO;
assign and_u1578_u0=and_u1576_u0&GO;
assign mux_u498=(and_u1577_u0)?add_u474:port_0002ea05_;
assign mux_u499_u0=(and_u1577_u0)?32'h0:add_u473;
assign simplePinWrite=reg_00b48d11_u0&{1{reg_00b48d11_u0}};
assign simplePinWrite_u237=port_00f9e1da_;
assign simplePinWrite_u238=16'h1&{16{1'h1}};
assign simplePinWrite_u239=16'h1&{16{1'h1}};
assign simplePinWrite_u240=port_0122d684_;
assign simplePinWrite_u241=reg_00b48d11_u0&{1{reg_00b48d11_u0}};
assign simplePinWrite_u242=reg_00b48d11_u0&{1{reg_00b48d11_u0}};
assign simplePinWrite_u243=16'h1&{16{1'h1}};
assign simplePinWrite_u244=port_002687bf_;
always @(posedge CLK)
begin
if (GO)
syncEnable_u360<=add_u464;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u361_u0<=add_u468;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00b48d11_u0<=1'h0;
else reg_00b48d11_u0<=reg_013422da_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_013422da_u0<=1'h0;
else reg_013422da_u0<=GO;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u362_u0<=add_u472;
end
assign RESULT=GO;
assign RESULT_u1006=mux_u498;
assign RESULT_u1007=GO;
assign RESULT_u1008=mux_u499_u0;
assign RESULT_u1009=reg_013422da_u0;
assign RESULT_u1010=syncEnable_u360;
assign RESULT_u1011=3'h1;
assign RESULT_u1012=reg_013422da_u0;
assign RESULT_u1013=syncEnable_u361_u0;
assign RESULT_u1014=3'h1;
assign RESULT_u1015=reg_013422da_u0;
assign RESULT_u1016=syncEnable_u362_u0;
assign RESULT_u1017=3'h1;
assign RESULT_u1018=simplePinWrite;
assign RESULT_u1019=simplePinWrite_u241;
assign RESULT_u1020=simplePinWrite_u244;
assign RESULT_u1021=simplePinWrite_u237;
assign RESULT_u1022=simplePinWrite_u243;
assign RESULT_u1023=simplePinWrite_u242;
assign RESULT_u1024=simplePinWrite_u238;
assign RESULT_u1025=simplePinWrite_u239;
assign RESULT_u1026=simplePinWrite_u240;
assign DONE=reg_00b48d11_u0;
endmodule



module output_process_Draw_rectangle_globalreset_physical_001fa2b7_(bus_0023db22_, bus_0113813a_, bus_00826511_);
input		bus_0023db22_;
input		bus_0113813a_;
output		bus_00826511_;
reg		sample_u21=1'h0;
wire		not_00f16943_u0;
reg		cross_u21=1'h0;
reg		final_u21=1'h1;
wire		and_0139d68e_u0;
reg		glitch_u21=1'h0;
wire		or_01890f98_u0;
always @(posedge bus_0023db22_)
begin
sample_u21<=1'h1;
end
assign bus_00826511_=or_01890f98_u0;
assign not_00f16943_u0=~and_0139d68e_u0;
always @(posedge bus_0023db22_)
begin
cross_u21<=sample_u21;
end
always @(posedge bus_0023db22_)
begin
final_u21<=not_00f16943_u0;
end
assign and_0139d68e_u0=cross_u21&glitch_u21;
always @(posedge bus_0023db22_)
begin
glitch_u21<=cross_u21;
end
assign or_01890f98_u0=bus_0113813a_|final_u21;
endmodule



module output_process_Draw_rectangle_drawRectangle(CLK, RESET, GO, port_00be099f_, port_0116e071_, port_000bb648_, port_01d67dc6_, port_01a2503a_, port_00891739_, port_0087f92c_, port_018e9e2f_, RESULT, RESULT_u1027, RESULT_u1028, RESULT_u1029, RESULT_u1030, RESULT_u1031, RESULT_u1032, RESULT_u1033, RESULT_u1034, RESULT_u1035, RESULT_u1036, RESULT_u1037, RESULT_u1038, RESULT_u1039, RESULT_u1040, RESULT_u1041, RESULT_u1042, RESULT_u1043, RESULT_u1044, RESULT_u1045, RESULT_u1046, RESULT_u1047, RESULT_u1048, RESULT_u1049, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_00be099f_;
input	[15:0]	port_0116e071_;
input		port_000bb648_;
input		port_01d67dc6_;
input		port_01a2503a_;
input		port_00891739_;
input		port_0087f92c_;
input		port_018e9e2f_;
output		RESULT;
output	[31:0]	RESULT_u1027;
output	[7:0]	RESULT_u1028;
output	[2:0]	RESULT_u1029;
output		RESULT_u1030;
output	[31:0]	RESULT_u1031;
output	[7:0]	RESULT_u1032;
output	[2:0]	RESULT_u1033;
output		RESULT_u1034;
output	[31:0]	RESULT_u1035;
output	[7:0]	RESULT_u1036;
output	[2:0]	RESULT_u1037;
output		RESULT_u1038;
output	[31:0]	RESULT_u1039;
output	[7:0]	RESULT_u1040;
output	[2:0]	RESULT_u1041;
output		RESULT_u1042;
output	[31:0]	RESULT_u1043;
output	[7:0]	RESULT_u1044;
output	[2:0]	RESULT_u1045;
output		RESULT_u1046;
output	[31:0]	RESULT_u1047;
output	[7:0]	RESULT_u1048;
output	[2:0]	RESULT_u1049;
output		DONE;
wire	[16:0]	subtract;
wire	[16:0]	subtract_u95;
wire	[16:0]	add;
wire	[16:0]	add_u475;
reg		reg_005dcf27_u0=1'h0;
reg		reg_005dcf27_result_delayed_u0=1'h0;
wire		and_u1579_u0;
wire	[31:0]	add_u476;
wire	[31:0]	add_u477;
wire	[31:0]	add_u478;
wire	[31:0]	add_u479;
wire		and_u1580_u0;
wire		or_u437_u0;
reg		reg_0137a99d_u0=1'h0;
wire	[31:0]	add_u480;
wire	[31:0]	add_u481;
wire	[31:0]	add_u482;
wire	[31:0]	add_u483;
wire		or_u438_u0;
wire		and_u1581_u0;
reg		reg_01cc78e9_u0=1'h0;
wire	[31:0]	add_u484;
wire	[31:0]	add_u485;
wire	[31:0]	add_u486;
wire	[31:0]	add_u487;
wire		and_u1582_u0;
wire		or_u439_u0;
reg		reg_019b6cf6_u0=1'h0;
wire	[31:0]	add_u488;
wire	[31:0]	add_u489;
wire	[31:0]	add_u490;
wire	[31:0]	add_u491;
wire		or_u440_u0;
reg		reg_01db7347_u0=1'h0;
wire		and_u1583_u0;
wire	[31:0]	add_u492;
wire	[31:0]	add_u493;
wire	[31:0]	add_u494;
wire	[31:0]	add_u495;
wire		and_u1584_u0;
wire		or_u441_u0;
reg		reg_01186c18_u0=1'h0;
wire	[31:0]	add_u496;
wire	[31:0]	add_u497;
wire	[31:0]	add_u498;
wire	[31:0]	add_u499;
reg		reg_00619e1f_u0=1'h0;
wire		or_u442_u0;
wire		and_u1585_u0;
wire	[31:0]	add_u500;
reg	[31:0]	syncEnable_u363=32'h0;
reg	[31:0]	syncEnable_u364_u0=32'h0;
reg		reg_01dddf42_u0=1'h0;
reg	[31:0]	syncEnable_u365_u0=32'h0;
reg	[31:0]	syncEnable_u366_u0=32'h0;
reg	[31:0]	syncEnable_u367_u0=32'h0;
reg	[31:0]	syncEnable_u368_u0=32'h0;
reg	[31:0]	syncEnable_u369_u0=32'h0;
reg		block_GO_delayed_u44=1'h0;
reg		and_delayed_u70=1'h0;
wire		and_u1586_u0;
wire signed	[31:0]	lessThanEqualTo_b_signed;
wire signed	[31:0]	lessThanEqualTo_a_signed;
wire		lessThanEqualTo;
wire		not_u326_u0;
wire		and_u1587_u0;
wire		and_u1588_u0;
reg	[17:0]	latch_007d61b9_reg=18'h0;
wire	[27:0]	latch_007d61b9_out;
wire	[31:0]	latch_001fc64b_out;
reg	[17:0]	latch_001fc64b_reg=18'h0;
reg	[16:0]	latch_00abd02d_reg=17'h0;
wire	[27:0]	latch_00abd02d_out;
wire		or_u443_u0;
wire	[31:0]	mux_u500;
reg		reg_0123d531_u0=1'h0;
reg		reg_012a167e_u0=1'h0;
wire	[31:0]	add_u501;
wire	[31:0]	add_u502;
wire	[31:0]	add_u503;
wire	[31:0]	add_u504;
wire		and_u1589_u0;
wire		or_u444_u0;
reg		reg_00aca92e_u0=1'h0;
wire	[31:0]	add_u505;
wire	[31:0]	add_u506;
wire	[31:0]	add_u507;
wire	[31:0]	add_u508;
wire		and_u1590_u0;
reg		reg_00ecb0f2_u0=1'h0;
wire		or_u445_u0;
wire	[31:0]	add_u509;
wire	[31:0]	add_u510;
wire	[31:0]	add_u511;
wire	[31:0]	add_u512;
wire		and_u1591_u0;
wire		or_u446_u0;
reg		reg_0098863f_u0=1'h0;
wire	[31:0]	add_u513;
wire	[31:0]	add_u514;
wire	[31:0]	add_u515;
wire	[31:0]	add_u516;
wire		and_u1592_u0;
wire		or_u447_u0;
reg		reg_01a5dc20_u0=1'h0;
wire	[31:0]	add_u517;
wire	[31:0]	add_u518;
wire	[31:0]	add_u519;
wire	[31:0]	add_u520;
wire		and_u1593_u0;
wire		or_u448_u0;
reg		reg_014b1a2e_u0=1'h0;
wire	[31:0]	add_u521;
wire	[31:0]	add_u522;
wire	[31:0]	add_u523;
wire	[31:0]	add_u524;
wire		or_u449_u0;
reg		reg_0112dff5_u0=1'h0;
wire		and_u1594_u0;
wire	[31:0]	add_u525;
reg	[31:0]	syncEnable_u370_u0=32'h0;
reg	[31:0]	syncEnable_u371_u0=32'h0;
reg		block_GO_delayed_u45_u0=1'h0;
reg	[31:0]	syncEnable_u372_u0=32'h0;
reg	[31:0]	syncEnable_u373_u0=32'h0;
reg		block_GO_delayed_result_delayed_u4=1'h0;
reg	[31:0]	syncEnable_u374_u0=32'h0;
reg	[31:0]	syncEnable_u375_u0=32'h0;
reg	[31:0]	syncEnable_u376_u0=32'h0;
wire		and_u1595_u0;
wire		lessThanEqualTo_u29;
wire signed	[31:0]	lessThanEqualTo_u29_b_signed;
wire signed	[31:0]	lessThanEqualTo_u29_a_signed;
wire		and_u1596_u0;
wire		and_u1597_u0;
wire		not_u327_u0;
reg		reg_012a167e_result_delayed_u0=1'h0;
wire		and_u1598_u0;
wire	[31:0]	latch_01348d26_out;
reg	[17:0]	latch_01348d26_reg=18'h0;
wire	[31:0]	latch_014ade69_out;
reg	[17:0]	latch_014ade69_reg=18'h0;
wire	[31:0]	latch_004cd203_out;
reg	[16:0]	latch_004cd203_reg=17'h0;
wire		or_u450_u0;
wire	[31:0]	mux_u501_u0;
reg	[17:0]	syncEnable_u377_u0=18'h0;
wire	[31:0]	mux_u502_u0;
wire		or_u451_u0;
wire	[31:0]	mux_u503_u0;
wire		or_u452_u0;
reg	[16:0]	syncEnable_u378_u0=17'h0;
wire		or_u453_u0;
wire	[31:0]	mux_u504_u0;
reg	[17:0]	syncEnable_u379_u0=18'h0;
reg		reg_0072cc7a_u0=1'h0;
wire	[31:0]	mux_u505_u0;
wire		or_u454_u0;
wire		or_u455_u0;
wire	[31:0]	mux_u506_u0;
wire	[31:0]	mux_u507_u0;
wire		or_u456_u0;
reg	[16:0]	syncEnable_u380_u0=17'h0;
assign subtract={1'b0, port_0116e071_}-17'ha;
assign subtract_u95={1'b0, port_00be099f_}-17'hd;
assign add={1'b0, port_0116e071_}+17'ha;
assign add_u475={1'b0, port_00be099f_}+17'hd;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_005dcf27_u0<=1'h0;
else reg_005dcf27_u0<=and_delayed_u70;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_005dcf27_result_delayed_u0<=1'h0;
else reg_005dcf27_result_delayed_u0<=reg_005dcf27_u0;
end
assign and_u1579_u0=and_u1587_u0&or_u443_u0;
assign add_u476={latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16:0], 7'b0}+{latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16:0], 5'b0};
assign add_u477={add_u476[24], add_u476[24], add_u476[24], add_u476[24], add_u476[24], add_u476[24], add_u476[24], add_u476[24:5], 5'b0}+{latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16:0], 4'b0};
assign add_u478={add_u477[25], add_u477[25], add_u477[25], add_u477[25], add_u477[25], add_u477[25], add_u477[25:4], 4'b0}+mux_u500;
assign add_u479=32'h0+add_u478;
assign and_u1580_u0=reg_0137a99d_u0&port_000bb648_;
assign or_u437_u0=and_u1580_u0|RESET;
always @(posedge CLK or posedge block_GO_delayed_u44 or posedge or_u437_u0)
begin
if (or_u437_u0)
reg_0137a99d_u0<=1'h0;
else if (block_GO_delayed_u44)
reg_0137a99d_u0<=1'h1;
else reg_0137a99d_u0<=reg_0137a99d_u0;
end
assign add_u480={latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16:0], 7'b0}+{latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16:0], 5'b0};
assign add_u481={add_u480[24], add_u480[24], add_u480[24], add_u480[24], add_u480[24], add_u480[24], add_u480[24], add_u480[24:5], 5'b0}+{latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16:0], 4'b0};
assign add_u482={add_u481[25], add_u481[25], add_u481[25], add_u481[25], add_u481[25], add_u481[25], add_u481[25:4], 4'b0}+mux_u500;
assign add_u483=32'h0+add_u482;
assign or_u438_u0=and_u1581_u0|RESET;
assign and_u1581_u0=reg_01cc78e9_u0&port_01d67dc6_;
always @(posedge CLK or posedge block_GO_delayed_u44 or posedge or_u438_u0)
begin
if (or_u438_u0)
reg_01cc78e9_u0<=1'h0;
else if (block_GO_delayed_u44)
reg_01cc78e9_u0<=1'h1;
else reg_01cc78e9_u0<=reg_01cc78e9_u0;
end
assign add_u484={latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16:0], 7'b0}+{latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16:0], 5'b0};
assign add_u485={add_u484[24], add_u484[24], add_u484[24], add_u484[24], add_u484[24], add_u484[24], add_u484[24], add_u484[24:5], 5'b0}+{latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16], latch_00abd02d_out[16:0], 4'b0};
assign add_u486={add_u485[25], add_u485[25], add_u485[25], add_u485[25], add_u485[25], add_u485[25], add_u485[25:4], 4'b0}+mux_u500;
assign add_u487=32'h0+add_u486;
assign and_u1582_u0=reg_019b6cf6_u0&port_01a2503a_;
assign or_u439_u0=and_u1582_u0|RESET;
always @(posedge CLK or posedge block_GO_delayed_u44 or posedge or_u439_u0)
begin
if (or_u439_u0)
reg_019b6cf6_u0<=1'h0;
else if (block_GO_delayed_u44)
reg_019b6cf6_u0<=1'h1;
else reg_019b6cf6_u0<=reg_019b6cf6_u0;
end
assign add_u488={8'b0, latch_007d61b9_out[16:0], 7'b0}+{10'b0, latch_007d61b9_out[16:0], 5'b0};
assign add_u489={add_u488[25], add_u488[25], add_u488[25], add_u488[25], add_u488[25], add_u488[25], add_u488[25:5], 5'b0}+{11'b0, latch_007d61b9_out[16:0], 4'b0};
assign add_u490={add_u489[26], add_u489[26], add_u489[26], add_u489[26], add_u489[26], add_u489[26:4], 4'b0}+mux_u500;
assign add_u491=32'h0+add_u490;
assign or_u440_u0=and_u1583_u0|RESET;
always @(posedge CLK or posedge reg_01dddf42_u0 or posedge or_u440_u0)
begin
if (or_u440_u0)
reg_01db7347_u0<=1'h0;
else if (reg_01dddf42_u0)
reg_01db7347_u0<=1'h1;
else reg_01db7347_u0<=reg_01db7347_u0;
end
assign and_u1583_u0=reg_01db7347_u0&port_00891739_;
assign add_u492={8'b0, latch_007d61b9_out[16:0], 7'b0}+{10'b0, latch_007d61b9_out[16:0], 5'b0};
assign add_u493={add_u492[25], add_u492[25], add_u492[25], add_u492[25], add_u492[25], add_u492[25], add_u492[25:5], 5'b0}+{11'b0, latch_007d61b9_out[16:0], 4'b0};
assign add_u494={add_u493[26], add_u493[26], add_u493[26], add_u493[26], add_u493[26], add_u493[26:4], 4'b0}+mux_u500;
assign add_u495=32'h0+add_u494;
assign and_u1584_u0=reg_01186c18_u0&port_018e9e2f_;
assign or_u441_u0=and_u1584_u0|RESET;
always @(posedge CLK or posedge reg_01dddf42_u0 or posedge or_u441_u0)
begin
if (or_u441_u0)
reg_01186c18_u0<=1'h0;
else if (reg_01dddf42_u0)
reg_01186c18_u0<=1'h1;
else reg_01186c18_u0<=reg_01186c18_u0;
end
assign add_u496={8'b0, latch_007d61b9_out[16:0], 7'b0}+{10'b0, latch_007d61b9_out[16:0], 5'b0};
assign add_u497={add_u496[25], add_u496[25], add_u496[25], add_u496[25], add_u496[25], add_u496[25], add_u496[25:5], 5'b0}+{11'b0, latch_007d61b9_out[16:0], 4'b0};
assign add_u498={add_u497[26], add_u497[26], add_u497[26], add_u497[26], add_u497[26], add_u497[26:4], 4'b0}+mux_u500;
assign add_u499=32'h0+add_u498;
always @(posedge CLK or posedge reg_01dddf42_u0 or posedge or_u442_u0)
begin
if (or_u442_u0)
reg_00619e1f_u0<=1'h0;
else if (reg_01dddf42_u0)
reg_00619e1f_u0<=1'h1;
else reg_00619e1f_u0<=reg_00619e1f_u0;
end
assign or_u442_u0=and_u1585_u0|RESET;
assign and_u1585_u0=reg_00619e1f_u0&port_0087f92c_;
assign add_u500=mux_u500+32'h1;
always @(posedge CLK)
begin
if (and_u1579_u0)
syncEnable_u363<=add_u499;
end
always @(posedge CLK)
begin
if (and_u1579_u0)
syncEnable_u364_u0<=add_u483;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01dddf42_u0<=1'h0;
else reg_01dddf42_u0<=block_GO_delayed_u44;
end
always @(posedge CLK)
begin
if (and_u1579_u0)
syncEnable_u365_u0<=add_u479;
end
always @(posedge CLK)
begin
if (and_u1579_u0)
syncEnable_u366_u0<=add_u491;
end
always @(posedge CLK)
begin
if (and_u1579_u0)
syncEnable_u367_u0<=add_u500;
end
always @(posedge CLK)
begin
if (and_u1579_u0)
syncEnable_u368_u0<=add_u487;
end
always @(posedge CLK)
begin
if (and_u1579_u0)
syncEnable_u369_u0<=add_u495;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u44<=1'h0;
else block_GO_delayed_u44<=and_u1579_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u70<=1'h0;
else and_delayed_u70<=and_u1579_u0;
end
assign and_u1586_u0=and_u1588_u0&or_u443_u0;
assign lessThanEqualTo_a_signed=mux_u500;
assign lessThanEqualTo_b_signed={15'b0, latch_001fc64b_out[16:0]};
assign lessThanEqualTo=lessThanEqualTo_a_signed<=lessThanEqualTo_b_signed;
assign not_u326_u0=~lessThanEqualTo;
assign and_u1587_u0=or_u443_u0&lessThanEqualTo;
assign and_u1588_u0=or_u443_u0&not_u326_u0;
always @(posedge CLK)
begin
if (reg_0072cc7a_u0)
latch_007d61b9_reg<={1'b0, syncEnable_u377_u0[16:0]};
end
assign latch_007d61b9_out=(reg_0072cc7a_u0)?{11'b0, syncEnable_u377_u0[16:0]}:{11'b0, latch_007d61b9_reg[16:0]};
assign latch_001fc64b_out=(reg_0072cc7a_u0)?{15'b0, syncEnable_u379_u0[16:0]}:{15'b0, latch_001fc64b_reg[16:0]};
always @(posedge CLK)
begin
if (reg_0072cc7a_u0)
latch_001fc64b_reg<={1'b0, syncEnable_u379_u0[16:0]};
end
always @(posedge CLK)
begin
if (reg_0072cc7a_u0)
latch_00abd02d_reg<=syncEnable_u378_u0;
end
assign latch_00abd02d_out=(reg_0072cc7a_u0)?{syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0}:{latch_00abd02d_reg[16], latch_00abd02d_reg[16], latch_00abd02d_reg[16], latch_00abd02d_reg[16], latch_00abd02d_reg[16], latch_00abd02d_reg[16], latch_00abd02d_reg[16], latch_00abd02d_reg[16], latch_00abd02d_reg[16], latch_00abd02d_reg[16], latch_00abd02d_reg[16], latch_00abd02d_reg};
assign or_u443_u0=reg_0072cc7a_u0|reg_005dcf27_result_delayed_u0;
assign mux_u500=(reg_0072cc7a_u0)?{syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0}:syncEnable_u367_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0123d531_u0<=1'h0;
else reg_0123d531_u0<=reg_012a167e_result_delayed_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_012a167e_u0<=1'h0;
else reg_012a167e_u0<=and_u1595_u0;
end
assign add_u501={mux_u501_u0[24:0], 7'b0}+{mux_u501_u0[26:0], 5'b0};
assign add_u502={add_u501[31:5], 5'b0}+{mux_u501_u0[27:0], 4'b0};
assign add_u503={add_u502[31:4], 4'b0}+{latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16:0]};
assign add_u504=32'h0+add_u503;
assign and_u1589_u0=reg_00aca92e_u0&port_000bb648_;
assign or_u444_u0=and_u1589_u0|RESET;
always @(posedge CLK or posedge block_GO_delayed_u45_u0 or posedge or_u444_u0)
begin
if (or_u444_u0)
reg_00aca92e_u0<=1'h0;
else if (block_GO_delayed_u45_u0)
reg_00aca92e_u0<=1'h1;
else reg_00aca92e_u0<=reg_00aca92e_u0;
end
assign add_u505={mux_u501_u0[24:0], 7'b0}+{mux_u501_u0[26:0], 5'b0};
assign add_u506={add_u505[31:5], 5'b0}+{mux_u501_u0[27:0], 4'b0};
assign add_u507={add_u506[31:4], 4'b0}+{latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16:0]};
assign add_u508=32'h0+add_u507;
assign and_u1590_u0=reg_00ecb0f2_u0&port_01d67dc6_;
always @(posedge CLK or posedge block_GO_delayed_u45_u0 or posedge or_u445_u0)
begin
if (or_u445_u0)
reg_00ecb0f2_u0<=1'h0;
else if (block_GO_delayed_u45_u0)
reg_00ecb0f2_u0<=1'h1;
else reg_00ecb0f2_u0<=reg_00ecb0f2_u0;
end
assign or_u445_u0=and_u1590_u0|RESET;
assign add_u509={mux_u501_u0[24:0], 7'b0}+{mux_u501_u0[26:0], 5'b0};
assign add_u510={add_u509[31:5], 5'b0}+{mux_u501_u0[27:0], 4'b0};
assign add_u511={add_u510[31:4], 4'b0}+{latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16], latch_004cd203_out[16:0]};
assign add_u512=32'h0+add_u511;
assign and_u1591_u0=reg_0098863f_u0&port_01a2503a_;
assign or_u446_u0=and_u1591_u0|RESET;
always @(posedge CLK or posedge block_GO_delayed_u45_u0 or posedge or_u446_u0)
begin
if (or_u446_u0)
reg_0098863f_u0<=1'h0;
else if (block_GO_delayed_u45_u0)
reg_0098863f_u0<=1'h1;
else reg_0098863f_u0<=reg_0098863f_u0;
end
assign add_u513={mux_u501_u0[24:0], 7'b0}+{mux_u501_u0[26:0], 5'b0};
assign add_u514={add_u513[31:5], 5'b0}+{mux_u501_u0[27:0], 4'b0};
assign add_u515={add_u514[31:4], 4'b0}+{15'b0, latch_014ade69_out[16:0]};
assign add_u516=32'h0+add_u515;
assign and_u1592_u0=reg_01a5dc20_u0&port_00891739_;
assign or_u447_u0=and_u1592_u0|RESET;
always @(posedge CLK or posedge block_GO_delayed_result_delayed_u4 or posedge or_u447_u0)
begin
if (or_u447_u0)
reg_01a5dc20_u0<=1'h0;
else if (block_GO_delayed_result_delayed_u4)
reg_01a5dc20_u0<=1'h1;
else reg_01a5dc20_u0<=reg_01a5dc20_u0;
end
assign add_u517={mux_u501_u0[24:0], 7'b0}+{mux_u501_u0[26:0], 5'b0};
assign add_u518={add_u517[31:5], 5'b0}+{mux_u501_u0[27:0], 4'b0};
assign add_u519={add_u518[31:4], 4'b0}+{15'b0, latch_014ade69_out[16:0]};
assign add_u520=32'h0+add_u519;
assign and_u1593_u0=reg_014b1a2e_u0&port_018e9e2f_;
assign or_u448_u0=and_u1593_u0|RESET;
always @(posedge CLK or posedge block_GO_delayed_result_delayed_u4 or posedge or_u448_u0)
begin
if (or_u448_u0)
reg_014b1a2e_u0<=1'h0;
else if (block_GO_delayed_result_delayed_u4)
reg_014b1a2e_u0<=1'h1;
else reg_014b1a2e_u0<=reg_014b1a2e_u0;
end
assign add_u521={mux_u501_u0[24:0], 7'b0}+{mux_u501_u0[26:0], 5'b0};
assign add_u522={add_u521[31:5], 5'b0}+{mux_u501_u0[27:0], 4'b0};
assign add_u523={add_u522[31:4], 4'b0}+{15'b0, latch_014ade69_out[16:0]};
assign add_u524=32'h0+add_u523;
assign or_u449_u0=and_u1594_u0|RESET;
always @(posedge CLK or posedge block_GO_delayed_result_delayed_u4 or posedge or_u449_u0)
begin
if (or_u449_u0)
reg_0112dff5_u0<=1'h0;
else if (block_GO_delayed_result_delayed_u4)
reg_0112dff5_u0<=1'h1;
else reg_0112dff5_u0<=reg_0112dff5_u0;
end
assign and_u1594_u0=reg_0112dff5_u0&port_0087f92c_;
assign add_u525=mux_u501_u0+32'h1;
always @(posedge CLK)
begin
if (and_u1595_u0)
syncEnable_u370_u0<=add_u520;
end
always @(posedge CLK)
begin
if (and_u1595_u0)
syncEnable_u371_u0<=add_u516;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u45_u0<=1'h0;
else block_GO_delayed_u45_u0<=and_u1595_u0;
end
always @(posedge CLK)
begin
if (and_u1595_u0)
syncEnable_u372_u0<=add_u504;
end
always @(posedge CLK)
begin
if (and_u1595_u0)
syncEnable_u373_u0<=add_u524;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_result_delayed_u4<=1'h0;
else block_GO_delayed_result_delayed_u4<=block_GO_delayed_u45_u0;
end
always @(posedge CLK)
begin
if (and_u1595_u0)
syncEnable_u374_u0<=add_u508;
end
always @(posedge CLK)
begin
if (and_u1595_u0)
syncEnable_u375_u0<=add_u512;
end
always @(posedge CLK)
begin
if (and_u1595_u0)
syncEnable_u376_u0<=add_u525;
end
assign and_u1595_u0=and_u1597_u0&or_u450_u0;
assign lessThanEqualTo_u29_a_signed=mux_u501_u0;
assign lessThanEqualTo_u29_b_signed={15'b0, latch_01348d26_out[16:0]};
assign lessThanEqualTo_u29=lessThanEqualTo_u29_a_signed<=lessThanEqualTo_u29_b_signed;
assign and_u1596_u0=or_u450_u0&not_u327_u0;
assign and_u1597_u0=or_u450_u0&lessThanEqualTo_u29;
assign not_u327_u0=~lessThanEqualTo_u29;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_012a167e_result_delayed_u0<=1'h0;
else reg_012a167e_result_delayed_u0<=reg_012a167e_u0;
end
assign and_u1598_u0=and_u1596_u0&or_u450_u0;
assign latch_01348d26_out=(and_u1586_u0)?{15'b0, syncEnable_u377_u0[16:0]}:{15'b0, latch_01348d26_reg[16:0]};
always @(posedge CLK)
begin
if (and_u1586_u0)
latch_01348d26_reg<={1'b0, syncEnable_u377_u0[16:0]};
end
assign latch_014ade69_out=(and_u1586_u0)?{15'b0, syncEnable_u379_u0[16:0]}:{15'b0, latch_014ade69_reg[16:0]};
always @(posedge CLK)
begin
if (and_u1586_u0)
latch_014ade69_reg<={1'b0, syncEnable_u379_u0[16:0]};
end
assign latch_004cd203_out=(and_u1586_u0)?{syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0[16], syncEnable_u380_u0}:{latch_004cd203_reg[16], latch_004cd203_reg[16], latch_004cd203_reg[16], latch_004cd203_reg[16], latch_004cd203_reg[16], latch_004cd203_reg[16], latch_004cd203_reg[16], latch_004cd203_reg[16], latch_004cd203_reg[16], latch_004cd203_reg[16], latch_004cd203_reg[16], latch_004cd203_reg[16], latch_004cd203_reg[16], latch_004cd203_reg[16], latch_004cd203_reg[16], latch_004cd203_reg};
always @(posedge CLK)
begin
if (and_u1586_u0)
latch_004cd203_reg<=syncEnable_u380_u0;
end
assign or_u450_u0=and_u1586_u0|reg_0123d531_u0;
assign mux_u501_u0=(and_u1586_u0)?{syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0[16], syncEnable_u378_u0}:syncEnable_u376_u0;
always @(posedge CLK)
begin
if (GO)
syncEnable_u377_u0<={1'b0, add_u475};
end
assign mux_u502_u0=(block_GO_delayed_u44)?syncEnable_u365_u0:syncEnable_u372_u0;
assign or_u451_u0=block_GO_delayed_u44|block_GO_delayed_u45_u0;
assign mux_u503_u0=(reg_01dddf42_u0)?syncEnable_u363:syncEnable_u373_u0;
assign or_u452_u0=reg_01dddf42_u0|block_GO_delayed_result_delayed_u4;
always @(posedge CLK)
begin
if (GO)
syncEnable_u378_u0<=subtract_u95;
end
assign or_u453_u0=block_GO_delayed_u44|block_GO_delayed_u45_u0;
assign mux_u504_u0=(block_GO_delayed_u44)?syncEnable_u368_u0:syncEnable_u375_u0;
always @(posedge CLK)
begin
if (GO)
syncEnable_u379_u0<={1'b0, add};
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0072cc7a_u0<=1'h0;
else reg_0072cc7a_u0<=GO;
end
assign mux_u505_u0=(reg_01dddf42_u0)?syncEnable_u366_u0:syncEnable_u371_u0;
assign or_u454_u0=reg_01dddf42_u0|block_GO_delayed_result_delayed_u4;
assign or_u455_u0=reg_01dddf42_u0|block_GO_delayed_result_delayed_u4;
assign mux_u506_u0=(reg_01dddf42_u0)?syncEnable_u369_u0:syncEnable_u370_u0;
assign mux_u507_u0=(block_GO_delayed_u44)?syncEnable_u364_u0:syncEnable_u374_u0;
assign or_u456_u0=block_GO_delayed_u44|block_GO_delayed_u45_u0;
always @(posedge CLK)
begin
if (GO)
syncEnable_u380_u0<=subtract;
end
assign RESULT=or_u451_u0;
assign RESULT_u1027=mux_u502_u0;
assign RESULT_u1028=8'hff;
assign RESULT_u1029=3'h1;
assign RESULT_u1030=or_u456_u0;
assign RESULT_u1031=mux_u507_u0;
assign RESULT_u1032=8'h0;
assign RESULT_u1033=3'h1;
assign RESULT_u1034=or_u453_u0;
assign RESULT_u1035=mux_u504_u0;
assign RESULT_u1036=8'h0;
assign RESULT_u1037=3'h1;
assign RESULT_u1038=or_u454_u0;
assign RESULT_u1039=mux_u505_u0;
assign RESULT_u1040=8'hff;
assign RESULT_u1041=3'h1;
assign RESULT_u1042=or_u452_u0;
assign RESULT_u1043=mux_u503_u0;
assign RESULT_u1044=8'h0;
assign RESULT_u1045=3'h1;
assign RESULT_u1046=or_u455_u0;
assign RESULT_u1047=mux_u506_u0;
assign RESULT_u1048=8'h0;
assign RESULT_u1049=3'h1;
assign DONE=and_u1598_u0;
endmodule



module output_process_Draw_rectangle_getValueRGB(CLK, RESET, GO, port_00c91e9e_, port_00c1d6b4_, port_00aa595c_, port_01e0f363_, port_006e1316_, port_016b104e_, port_00a96b61_, port_004f15e5_, RESULT, RESULT_u1050, RESULT_u1051, RESULT_u1052, RESULT_u1053, RESULT_u1054, RESULT_u1055, RESULT_u1056, RESULT_u1057, RESULT_u1058, RESULT_u1059, RESULT_u1060, RESULT_u1061, RESULT_u1062, RESULT_u1063, RESULT_u1064, RESULT_u1065, RESULT_u1066, RESULT_u1067, DONE);
input		CLK;
input		RESET;
input		GO;
input	[31:0]	port_00c91e9e_;
input	[31:0]	port_00c1d6b4_;
input		port_00aa595c_;
input		port_01e0f363_;
input		port_006e1316_;
input	[7:0]	port_016b104e_;
input	[7:0]	port_00a96b61_;
input	[7:0]	port_004f15e5_;
output		RESULT;
output	[31:0]	RESULT_u1050;
output		RESULT_u1051;
output	[31:0]	RESULT_u1052;
output		RESULT_u1053;
output	[31:0]	RESULT_u1054;
output	[7:0]	RESULT_u1055;
output	[2:0]	RESULT_u1056;
output		RESULT_u1057;
output	[31:0]	RESULT_u1058;
output	[7:0]	RESULT_u1059;
output	[2:0]	RESULT_u1060;
output		RESULT_u1061;
output	[31:0]	RESULT_u1062;
output	[7:0]	RESULT_u1063;
output	[2:0]	RESULT_u1064;
output		RESULT_u1065;
output		RESULT_u1066;
output		RESULT_u1067;
output		DONE;
wire		simplePinWrite;
wire		simplePinWrite_u245;
wire		simplePinWrite_u246;
wire	[31:0]	add;
wire	[31:0]	add_u526;
wire	[31:0]	add_u527;
wire	[31:0]	add_u528;
wire		or_u457_u0;
wire		and_u1599_u0;
reg		reg_00bc8f4a_u0=1'h0;
wire	[31:0]	add_u529;
wire	[31:0]	add_u530;
wire	[31:0]	add_u531;
wire	[31:0]	add_u532;
wire		and_u1600_u0;
wire		or_u458_u0;
reg		reg_01f9ed0b_u0=1'h0;
wire	[31:0]	add_u533;
wire	[31:0]	add_u534;
wire	[31:0]	add_u535;
wire	[31:0]	add_u536;
wire		or_u459_u0;
wire		and_u1601_u0;
reg		reg_001b3cf1_u0=1'h0;
wire	[31:0]	add_u537;
wire signed	[31:0]	equals_b_signed;
wire signed	[31:0]	equals_a_signed;
wire		equals;
wire		and_u1602_u0;
wire		not_u328_u0;
wire		and_u1603_u0;
wire	[31:0]	add_u538;
wire	[31:0]	mux_u508;
wire		and_u1604_u0;
wire		and_u1605_u0;
wire	[31:0]	mux_u509_u0;
reg	[31:0]	syncEnable_u381=32'h0;
reg	[7:0]	syncEnable_u382_u0=8'h0;
reg		reg_018de1e2_u0=1'h0;
reg	[31:0]	syncEnable_u383_u0=32'h0;
reg	[7:0]	syncEnable_u384_u0=8'h0;
reg	[31:0]	syncEnable_u385_u0=32'h0;
reg		reg_01d915c1_u0=1'h0;
reg	[7:0]	syncEnable_u386_u0=8'h0;
assign simplePinWrite=GO&{1{GO}};
assign simplePinWrite_u245=GO&{1{GO}};
assign simplePinWrite_u246=GO&{1{GO}};
assign add={port_00c91e9e_[24:0], 7'b0}+{port_00c91e9e_[26:0], 5'b0};
assign add_u526={add[31:5], 5'b0}+{port_00c91e9e_[27:0], 4'b0};
assign add_u527={add_u526[31:4], 4'b0}+port_00c1d6b4_;
assign add_u528=32'h0+add_u527;
assign or_u457_u0=and_u1599_u0|RESET;
assign and_u1599_u0=reg_00bc8f4a_u0&port_00aa595c_;
always @(posedge CLK or posedge reg_01d915c1_u0 or posedge or_u457_u0)
begin
if (or_u457_u0)
reg_00bc8f4a_u0<=1'h0;
else if (reg_01d915c1_u0)
reg_00bc8f4a_u0<=1'h1;
else reg_00bc8f4a_u0<=reg_00bc8f4a_u0;
end
assign add_u529={port_00c91e9e_[24:0], 7'b0}+{port_00c91e9e_[26:0], 5'b0};
assign add_u530={add_u529[31:5], 5'b0}+{port_00c91e9e_[27:0], 4'b0};
assign add_u531={add_u530[31:4], 4'b0}+port_00c1d6b4_;
assign add_u532=32'h0+add_u531;
assign and_u1600_u0=reg_01f9ed0b_u0&port_01e0f363_;
assign or_u458_u0=and_u1600_u0|RESET;
always @(posedge CLK or posedge reg_01d915c1_u0 or posedge or_u458_u0)
begin
if (or_u458_u0)
reg_01f9ed0b_u0<=1'h0;
else if (reg_01d915c1_u0)
reg_01f9ed0b_u0<=1'h1;
else reg_01f9ed0b_u0<=reg_01f9ed0b_u0;
end
assign add_u533={port_00c91e9e_[24:0], 7'b0}+{port_00c91e9e_[26:0], 5'b0};
assign add_u534={add_u533[31:5], 5'b0}+{port_00c91e9e_[27:0], 4'b0};
assign add_u535={add_u534[31:4], 4'b0}+port_00c1d6b4_;
assign add_u536=32'h0+add_u535;
assign or_u459_u0=and_u1601_u0|RESET;
assign and_u1601_u0=reg_001b3cf1_u0&port_006e1316_;
always @(posedge CLK or posedge reg_01d915c1_u0 or posedge or_u459_u0)
begin
if (or_u459_u0)
reg_001b3cf1_u0<=1'h0;
else if (reg_01d915c1_u0)
reg_001b3cf1_u0<=1'h1;
else reg_001b3cf1_u0<=reg_001b3cf1_u0;
end
assign add_u537=port_00c1d6b4_+32'h1;
assign equals_a_signed=add_u537;
assign equals_b_signed=32'hb0;
assign equals=equals_a_signed==equals_b_signed;
assign and_u1602_u0=GO&not_u328_u0;
assign not_u328_u0=~equals;
assign and_u1603_u0=GO&equals;
assign add_u538=port_00c91e9e_+32'h1;
assign mux_u508=(and_u1604_u0)?port_00c91e9e_:add_u538;
assign and_u1604_u0=and_u1602_u0&GO;
assign and_u1605_u0=and_u1603_u0&GO;
assign mux_u509_u0=(and_u1604_u0)?add_u537:32'h0;
always @(posedge CLK)
begin
if (GO)
syncEnable_u381<=add_u532;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u382_u0<=port_016b104e_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_018de1e2_u0<=1'h0;
else reg_018de1e2_u0<=reg_01d915c1_u0;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u383_u0<=add_u528;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u384_u0<=port_004f15e5_;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u385_u0<=add_u536;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01d915c1_u0<=1'h0;
else reg_01d915c1_u0<=GO;
end
always @(posedge CLK)
begin
if (GO)
syncEnable_u386_u0<=port_00a96b61_;
end
assign RESULT=GO;
assign RESULT_u1050=mux_u508;
assign RESULT_u1051=GO;
assign RESULT_u1052=mux_u509_u0;
assign RESULT_u1053=reg_01d915c1_u0;
assign RESULT_u1054=syncEnable_u383_u0;
assign RESULT_u1055=syncEnable_u386_u0;
assign RESULT_u1056=3'h1;
assign RESULT_u1057=reg_01d915c1_u0;
assign RESULT_u1058=syncEnable_u381;
assign RESULT_u1059=syncEnable_u384_u0;
assign RESULT_u1060=3'h1;
assign RESULT_u1061=reg_01d915c1_u0;
assign RESULT_u1062=syncEnable_u385_u0;
assign RESULT_u1063=syncEnable_u382_u0;
assign RESULT_u1064=3'h1;
assign RESULT_u1065=simplePinWrite_u246;
assign RESULT_u1066=simplePinWrite_u245;
assign RESULT_u1067=simplePinWrite;
assign DONE=reg_018de1e2_u0;
endmodule



module output_process_Draw_rectangle_Kicker_21(CLK, RESET, bus_00e9d5a0_);
input		CLK;
input		RESET;
output		bus_00e9d5a0_;
wire		bus_01575c46_;
wire		bus_01118bc6_;
reg		kicker_2=1'h0;
wire		bus_003075b4_;
reg		kicker_res=1'h0;
reg		kicker_1=1'h0;
wire		bus_00dab253_;
assign bus_01575c46_=bus_00dab253_&kicker_1;
assign bus_01118bc6_=kicker_1&bus_00dab253_&bus_003075b4_;
always @(posedge CLK)
begin
kicker_2<=bus_01575c46_;
end
assign bus_00e9d5a0_=kicker_res;
assign bus_003075b4_=~kicker_2;
always @(posedge CLK)
begin
kicker_res<=bus_01118bc6_;
end
always @(posedge CLK)
begin
kicker_1<=bus_00dab253_;
end
assign bus_00dab253_=~RESET;
endmodule



module output_process_Draw_rectangle_simplememoryreferee_01bc888a_(bus_00150c03_, bus_01c7b9d3_, bus_01179579_, bus_01764864_, bus_00a40f07_, bus_00bb1f5c_, bus_010d3878_, bus_002943c5_, bus_008abdc8_, bus_015653dd_, bus_00c3bb80_, bus_00e4d935_, bus_014758cb_, bus_01203b9e_);
input		bus_00150c03_;
input		bus_01c7b9d3_;
input		bus_01179579_;
input	[7:0]	bus_01764864_;
input		bus_00a40f07_;
input	[7:0]	bus_00bb1f5c_;
input	[31:0]	bus_010d3878_;
input	[2:0]	bus_002943c5_;
output	[7:0]	bus_008abdc8_;
output	[31:0]	bus_015653dd_;
output		bus_00c3bb80_;
output		bus_00e4d935_;
output	[2:0]	bus_014758cb_;
output		bus_01203b9e_;
assign bus_008abdc8_=8'h0;
assign bus_015653dd_=bus_010d3878_;
assign bus_00c3bb80_=bus_00a40f07_;
assign bus_00e4d935_=bus_00a40f07_;
assign bus_014758cb_=3'h1;
assign bus_01203b9e_=bus_01179579_;
endmodule



module output_process_Draw_rectangle_structuralmemory_0198cbd9_(CLK_u42, bus_01d301f6_, bus_01c3d072_, bus_014da5cc_, bus_0169c6de_, bus_014ecd16_, bus_01437b60_, bus_01e5c110_, bus_00c30c8e_, bus_0143d8b1_, bus_0031ac17_, bus_017f3e79_, bus_015914b1_, bus_0119517f_);
input		CLK_u42;
input		bus_01d301f6_;
input	[31:0]	bus_01c3d072_;
input	[2:0]	bus_014da5cc_;
input		bus_0169c6de_;
input		bus_014ecd16_;
input	[7:0]	bus_01437b60_;
input	[31:0]	bus_01e5c110_;
input	[2:0]	bus_00c30c8e_;
input		bus_0143d8b1_;
input	[7:0]	bus_0031ac17_;
output	[7:0]	bus_017f3e79_;
output		bus_015914b1_;
output		bus_0119517f_;
reg		logicalMem_bbd522_we_delay0_u0=1'h0;
wire	[7:0]	bus_00bee7d6_;
wire		or_00828f12_u0;
reg		logicalMem_bbd522_re_delay0_u0=1'h0;
wire		or_01e2e881_u0;
reg		logicalMem_bbd522_we_delay0_u1_u0=1'h0;
always @(posedge CLK_u42 or posedge bus_01d301f6_)
begin
if (bus_01d301f6_)
logicalMem_bbd522_we_delay0_u0<=1'h0;
else logicalMem_bbd522_we_delay0_u0<=bus_0143d8b1_;
end
output_process_Draw_rectangle_forge_memory_25344x8_69 output_process_Draw_rectangle_forge_memory_25344x8_69_instance2(.CLK(CLK_u42), 
  .ENA(or_00828f12_u0), .WEA(bus_014ecd16_), .DINA(bus_01437b60_), .ADDRA(bus_01c3d072_), 
  .DOUTA(bus_00bee7d6_), .DONEA(), .ENB(bus_0143d8b1_), .WEB(bus_0143d8b1_), .DINB(8'hff), 
  .ADDRB(bus_01e5c110_), .DONEB());
assign or_00828f12_u0=bus_0169c6de_|bus_014ecd16_;
assign bus_017f3e79_=bus_00bee7d6_;
assign bus_015914b1_=or_01e2e881_u0;
assign bus_0119517f_=logicalMem_bbd522_we_delay0_u0;
always @(posedge CLK_u42 or posedge bus_01d301f6_)
begin
if (bus_01d301f6_)
logicalMem_bbd522_re_delay0_u0<=1'h0;
else logicalMem_bbd522_re_delay0_u0<=bus_0169c6de_;
end
assign or_01e2e881_u0=logicalMem_bbd522_re_delay0_u0|logicalMem_bbd522_we_delay0_u1_u0;
always @(posedge CLK_u42 or posedge bus_01d301f6_)
begin
if (bus_01d301f6_)
logicalMem_bbd522_we_delay0_u1_u0<=1'h0;
else logicalMem_bbd522_we_delay0_u1_u0<=bus_014ecd16_;
end
endmodule



module output_process_Draw_rectangle_endianswapper_00c13abb_(endianswapper_00c13abb_in, endianswapper_00c13abb_out);
input	[15:0]	endianswapper_00c13abb_in;
output	[15:0]	endianswapper_00c13abb_out;
assign endianswapper_00c13abb_out=endianswapper_00c13abb_in;
endmodule



module output_process_Draw_rectangle_endianswapper_00792464_(endianswapper_00792464_in, endianswapper_00792464_out);
input	[15:0]	endianswapper_00792464_in;
output	[15:0]	endianswapper_00792464_out;
assign endianswapper_00792464_out=endianswapper_00792464_in;
endmodule



module output_process_Draw_rectangle_stateVar_centre_y(bus_008068bf_, bus_005cd3da_, bus_002324b9_, bus_00e92383_, bus_01915a27_);
input		bus_008068bf_;
input		bus_005cd3da_;
input		bus_002324b9_;
input	[15:0]	bus_00e92383_;
output	[15:0]	bus_01915a27_;
wire	[15:0]	endianswapper_00c13abb_out;
reg	[15:0]	stateVar_centre_y_u5=16'h0;
wire	[15:0]	endianswapper_00792464_out;
assign bus_01915a27_=endianswapper_00792464_out;
output_process_Draw_rectangle_endianswapper_00c13abb_ output_process_Draw_rectangle_endianswapper_00c13abb__1(.endianswapper_00c13abb_in(bus_00e92383_), 
  .endianswapper_00c13abb_out(endianswapper_00c13abb_out));
always @(posedge bus_008068bf_ or posedge bus_005cd3da_)
begin
if (bus_005cd3da_)
stateVar_centre_y_u5<=16'h0;
else if (bus_002324b9_)
stateVar_centre_y_u5<=endianswapper_00c13abb_out;
end
output_process_Draw_rectangle_endianswapper_00792464_ output_process_Draw_rectangle_endianswapper_00792464__1(.endianswapper_00792464_in(stateVar_centre_y_u5), 
  .endianswapper_00792464_out(endianswapper_00792464_out));
endmodule



module output_process_Draw_rectangle_stateVar_state_s0(bus_012cd072_, bus_01290bbe_, bus_00c0ada5_, bus_002ce97c_, bus_0074d452_);
input		bus_012cd072_;
input		bus_01290bbe_;
input		bus_00c0ada5_;
input		bus_002ce97c_;
output		bus_0074d452_;
reg		stateVar_state_s0_u16=1'h0;
assign bus_0074d452_=stateVar_state_s0_u16;
always @(posedge bus_012cd072_ or posedge bus_01290bbe_)
begin
if (bus_01290bbe_)
stateVar_state_s0_u16<=1'h0;
else if (bus_00c0ada5_)
stateVar_state_s0_u16<=bus_002ce97c_;
end
endmodule



module output_process_Draw_rectangle_simplememoryreferee_00d7a4d7_(bus_0121612e_, bus_00732c35_, bus_009da5d7_, bus_005076d2_, bus_0188d17c_, bus_0138f3bb_, bus_01d679a0_, bus_00aa30fc_, bus_00a8f1e0_, bus_00b4f835_, bus_01ff134d_, bus_008cf4be_, bus_0076b457_, bus_0176022b_);
input		bus_0121612e_;
input		bus_00732c35_;
input		bus_009da5d7_;
input	[7:0]	bus_005076d2_;
input		bus_0188d17c_;
input	[7:0]	bus_0138f3bb_;
input	[31:0]	bus_01d679a0_;
input	[2:0]	bus_00aa30fc_;
output	[7:0]	bus_00a8f1e0_;
output	[31:0]	bus_00b4f835_;
output		bus_01ff134d_;
output		bus_008cf4be_;
output	[2:0]	bus_0076b457_;
output		bus_0176022b_;
assign bus_00a8f1e0_=8'h0;
assign bus_00b4f835_=bus_01d679a0_;
assign bus_01ff134d_=bus_0188d17c_;
assign bus_008cf4be_=bus_0188d17c_;
assign bus_0076b457_=3'h1;
assign bus_0176022b_=bus_009da5d7_;
endmodule



module output_process_Draw_rectangle_stateVar_state_s2(bus_00f238fa_, bus_007ac458_, bus_005d6340_, bus_000dff53_, bus_01cd028e_);
input		bus_00f238fa_;
input		bus_007ac458_;
input		bus_005d6340_;
input		bus_000dff53_;
output		bus_01cd028e_;
reg		stateVar_state_s2_u10=1'h0;
assign bus_01cd028e_=stateVar_state_s2_u10;
always @(posedge bus_00f238fa_ or posedge bus_007ac458_)
begin
if (bus_007ac458_)
stateVar_state_s2_u10<=1'h0;
else if (bus_005d6340_)
stateVar_state_s2_u10<=bus_000dff53_;
end
endmodule



module output_process_Draw_rectangle_scheduler(CLK, RESET, GO, port_003e9bda_, port_01961eea_, port_0012bfe7_, port_0055998f_, port_01f67390_, port_000bbff8_, port_01b61592_, port_0091ced8_, port_002e8e34_, port_01613518_, port_0192ec25_, port_01ca5227_, port_01559388_, port_00cb09f8_, port_01572c5f_, port_012d89fe_, port_009db78a_, port_007e9851_, RESULT, RESULT_u1068, RESULT_u1069, RESULT_u1070, RESULT_u1071, RESULT_u1072, RESULT_u1073, RESULT_u1074, RESULT_u1075, RESULT_u1076, RESULT_u1077, RESULT_u1078, RESULT_u1079, DONE);
input		CLK;
input		RESET;
input		GO;
input		port_003e9bda_;
input		port_01961eea_;
input		port_0012bfe7_;
input		port_0055998f_;
input	[31:0]	port_01f67390_;
input		port_000bbff8_;
input		port_01b61592_;
input		port_0091ced8_;
input		port_002e8e34_;
input		port_01613518_;
input		port_0192ec25_;
input		port_01ca5227_;
input		port_01559388_;
input		port_00cb09f8_;
input		port_01572c5f_;
input		port_012d89fe_;
input		port_009db78a_;
input		port_007e9851_;
output		RESULT;
output		RESULT_u1068;
output		RESULT_u1069;
output		RESULT_u1070;
output		RESULT_u1071;
output		RESULT_u1072;
output		RESULT_u1073;
output		RESULT_u1074;
output		RESULT_u1075;
output		RESULT_u1076;
output		RESULT_u1077;
output		RESULT_u1078;
output		RESULT_u1079;
output		DONE;
wire		and_u1606_u0;
wire		and_u1607_u0;
wire		and_u1608_u0;
wire		and_u1609_u0;
wire signed	[31:0]	equals_b_signed;
wire signed	[31:0]	equals_a_signed;
wire		equals;
wire		and_u1610_u0;
wire		and_u1611_u0;
wire		and_u1612_u0;
wire		and_u1613_u0;
wire		not_u329_u0;
wire		and_u1614_u0;
wire		not_u330_u0;
wire		and_u1615_u0;
wire		simplePinWrite;
wire		and_u1616_u0;
wire		and_u1617_u0;
wire		not_u331_u0;
wire		and_u1618_u0;
wire		simplePinWrite_u247;
wire		and_u1619_u0;
wire		or_u460_u0;
wire		and_u1620_u0;
reg		reg_0036baae_u0=1'h0;
reg		reg_00921baf_u0=1'h0;
reg		and_delayed_u71=1'h0;
wire		and_u1621_u0;
wire		and_u1622_u0;
wire		or_u461_u0;
reg		and_delayed_u72_u0=1'h0;
wire		and_u1623_u0;
reg		reg_00dc96b7_u0=1'h0;
wire		and_u1624_u0;
wire		and_u1625_u0;
wire		or_u462_u0;
wire		and_u1626_u0;
wire		and_u1627_u0;
wire		not_u332_u0;
wire		and_u1628_u0;
wire		not_u333_u0;
wire		and_u1629_u0;
wire		simplePinWrite_u248;
wire		and_u1630_u0;
wire		and_u1631_u0;
wire		and_u1632_u0;
wire		and_u1633_u0;
wire		not_u334_u0;
wire		and_u1634_u0;
wire		simplePinWrite_u249;
wire		and_u1635_u0;
wire		and_u1636_u0;
wire		and_u1637_u0;
reg		reg_00a4a314_u0=1'h0;
wire		and_u1638_u0;
wire		or_u463_u0;
wire		not_u335_u0;
wire		and_u1639_u0;
wire		and_u1640_u0;
wire		not_u336_u0;
wire		and_u1641_u0;
wire		and_u1642_u0;
wire		simplePinWrite_u250;
wire		and_u1643_u0;
wire		and_u1644_u0;
wire		and_u1645_u0;
wire		not_u337_u0;
wire		simplePinWrite_u251;
reg		reg_012b2be0_u0=1'h0;
reg		reg_01df33da_u0=1'h0;
wire		or_u464_u0;
wire		and_u1646_u0;
wire		and_u1647_u0;
reg		reg_012b2be0_result_delayed_u0=1'h0;
wire		and_u1648_u0;
wire		or_u465_u0;
wire		and_u1649_u0;
reg		reg_00040e54_u0=1'h0;
wire		and_u1650_u0;
reg		reg_012e842a_u0=1'h0;
wire		and_u1651_u0;
wire		and_u1652_u0;
wire		or_u466_u0;
wire		scoreboard_00157922_resOr2;
wire		scoreboard_00157922_resOr0;
reg		scoreboard_00157922_reg2=1'h0;
reg		scoreboard_00157922_reg1=1'h0;
wire		scoreboard_00157922_and;
wire		bus_001fcb73_;
wire		scoreboard_00157922_resOr1;
reg		scoreboard_00157922_reg0=1'h0;
wire		doneCountIm_go_merge;
wire		mux_u510;
wire		or_u467_u0;
wire		or_u468_u0;
wire		mux_u511_u0;
wire		or_u469_u0;
wire		mux_u512_u0;
wire		or_u470_u0;
wire		mux_u513_u0;
reg		syncEnable_u387=1'h0;
reg		syncEnable_u388_u0=1'h0;
reg		syncEnable_u389_u0=1'h0;
reg		syncEnable_u390_u0=1'h0;
reg		syncEnable_u391_u0=1'h0;
reg		syncEnable_u392_u0=1'h0;
reg		block_GO_delayed_u46=1'h0;
reg		syncEnable_u393_u0=1'h0;
reg		syncEnable_u394_u0=1'h0;
wire		or_u471_u0;
reg		loopControl_u35=1'h0;
wire		or_u472_u0;
wire		mux_u514_u0;
reg		reg_0122bb99_u0=1'h0;
wire		or_u473_u0;
wire		mux_u515_u0;
reg		reg_006b4712_u0=1'h0;
wire		or_u474_u0;
wire		mux_u516_u0;
wire		or_u475_u0;
wire		mux_u517_u0;
assign and_u1606_u0=or_u471_u0&or_u471_u0;
assign and_u1607_u0=port_000bbff8_&port_01ca5227_;
assign and_u1608_u0=port_002e8e34_&port_0192ec25_;
assign and_u1609_u0=and_u1608_u0&port_01613518_;
assign equals_a_signed=port_01f67390_;
assign equals_b_signed=32'h90;
assign equals=equals_a_signed==equals_b_signed;
assign and_u1610_u0=port_01559388_&port_01572c5f_;
assign and_u1611_u0=and_u1610_u0&port_009db78a_;
assign and_u1612_u0=block_GO_delayed_u46&not_u329_u0;
assign and_u1613_u0=block_GO_delayed_u46&syncEnable_u387;
assign not_u329_u0=~syncEnable_u387;
assign and_u1614_u0=and_u1624_u0&not_u330_u0;
assign not_u330_u0=~syncEnable_u393_u0;
assign and_u1615_u0=and_u1624_u0&syncEnable_u393_u0;
assign simplePinWrite=and_u1616_u0&{1{and_u1616_u0}};
assign and_u1616_u0=and_u1622_u0&and_u1622_u0;
assign and_u1617_u0=and_u1623_u0&not_u331_u0;
assign not_u331_u0=~syncEnable_u390_u0;
assign and_u1618_u0=and_u1623_u0&syncEnable_u390_u0;
assign simplePinWrite_u247=and_u1619_u0&{1{and_u1619_u0}};
assign and_u1619_u0=and_u1621_u0&and_u1621_u0;
assign or_u460_u0=and_delayed_u71|reg_0036baae_u0;
assign and_u1620_u0=and_u1617_u0&and_u1623_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0036baae_u0<=1'h0;
else reg_0036baae_u0<=reg_00921baf_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00921baf_u0<=1'h0;
else reg_00921baf_u0<=and_u1621_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u71<=1'h0;
else and_delayed_u71<=and_u1620_u0;
end
assign and_u1621_u0=and_u1618_u0&and_u1623_u0;
assign and_u1622_u0=and_u1615_u0&and_u1624_u0;
assign or_u461_u0=or_u460_u0|and_delayed_u72_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
and_delayed_u72_u0<=1'h0;
else and_delayed_u72_u0<=and_u1622_u0;
end
assign and_u1623_u0=and_u1614_u0&and_u1624_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00dc96b7_u0<=1'h0;
else reg_00dc96b7_u0<=and_u1625_u0;
end
assign and_u1624_u0=and_u1613_u0&block_GO_delayed_u46;
assign and_u1625_u0=and_u1612_u0&block_GO_delayed_u46;
assign or_u462_u0=or_u461_u0|reg_00dc96b7_u0;
assign and_u1626_u0=block_GO_delayed_u46&not_u332_u0;
assign and_u1627_u0=block_GO_delayed_u46&syncEnable_u389_u0;
assign not_u332_u0=~syncEnable_u389_u0;
assign and_u1628_u0=and_u1632_u0&not_u333_u0;
assign not_u333_u0=~syncEnable_u388_u0;
assign and_u1629_u0=and_u1632_u0&syncEnable_u388_u0;
assign simplePinWrite_u248=and_u1630_u0&{1{and_u1630_u0}};
assign and_u1630_u0=and_u1631_u0&and_u1631_u0;
assign and_u1631_u0=and_u1629_u0&and_u1632_u0;
assign and_u1632_u0=and_u1627_u0&block_GO_delayed_u46;
assign and_u1633_u0=block_GO_delayed_u46&not_u334_u0;
assign not_u334_u0=~syncEnable_u392_u0;
assign and_u1634_u0=block_GO_delayed_u46&syncEnable_u392_u0;
assign simplePinWrite_u249=and_u1635_u0&{1{and_u1635_u0}};
assign and_u1635_u0=and_u1636_u0&and_u1636_u0;
assign and_u1636_u0=and_u1637_u0&and_u1637_u0;
assign and_u1637_u0=and_u1634_u0&block_GO_delayed_u46;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00a4a314_u0<=1'h0;
else reg_00a4a314_u0<=and_u1638_u0;
end
assign and_u1638_u0=and_u1633_u0&block_GO_delayed_u46;
assign or_u463_u0=port_012d89fe_|reg_00a4a314_u0;
assign not_u335_u0=~syncEnable_u391_u0;
assign and_u1639_u0=block_GO_delayed_u46&not_u335_u0;
assign and_u1640_u0=block_GO_delayed_u46&syncEnable_u391_u0;
assign not_u336_u0=~syncEnable_u393_u0;
assign and_u1641_u0=and_u1651_u0&not_u336_u0;
assign and_u1642_u0=and_u1651_u0&syncEnable_u393_u0;
assign simplePinWrite_u250=and_u1643_u0&{1{and_u1643_u0}};
assign and_u1643_u0=and_u1650_u0&and_u1650_u0;
assign and_u1644_u0=and_u1648_u0&not_u337_u0;
assign and_u1645_u0=and_u1648_u0&and_u1611_u0;
assign not_u337_u0=~and_u1611_u0;
assign simplePinWrite_u251=and_u1646_u0&{1{and_u1646_u0}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_012b2be0_u0<=1'h0;
else reg_012b2be0_u0<=and_u1646_u0;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_01df33da_u0<=1'h0;
else reg_01df33da_u0<=and_u1647_u0;
end
assign or_u464_u0=reg_012b2be0_result_delayed_u0|reg_01df33da_u0;
assign and_u1646_u0=and_u1645_u0&and_u1648_u0;
assign and_u1647_u0=and_u1644_u0&and_u1648_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_012b2be0_result_delayed_u0<=1'h0;
else reg_012b2be0_result_delayed_u0<=reg_012b2be0_u0;
end
assign and_u1648_u0=and_u1649_u0&and_u1649_u0;
assign or_u465_u0=reg_00040e54_u0|or_u464_u0;
assign and_u1649_u0=and_u1641_u0&and_u1651_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00040e54_u0<=1'h0;
else reg_00040e54_u0<=and_u1650_u0;
end
assign and_u1650_u0=and_u1642_u0&and_u1651_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_012e842a_u0<=1'h0;
else reg_012e842a_u0<=and_u1652_u0;
end
assign and_u1651_u0=and_u1640_u0&block_GO_delayed_u46;
assign and_u1652_u0=and_u1639_u0&block_GO_delayed_u46;
assign or_u466_u0=or_u465_u0|reg_012e842a_u0;
assign scoreboard_00157922_resOr2=or_u463_u0|scoreboard_00157922_reg2;
assign scoreboard_00157922_resOr0=or_u466_u0|scoreboard_00157922_reg0;
always @(posedge CLK)
begin
if (bus_001fcb73_)
scoreboard_00157922_reg2<=1'h0;
else if (or_u463_u0)
scoreboard_00157922_reg2<=1'h1;
else scoreboard_00157922_reg2<=scoreboard_00157922_reg2;
end
always @(posedge CLK)
begin
if (bus_001fcb73_)
scoreboard_00157922_reg1<=1'h0;
else if (or_u462_u0)
scoreboard_00157922_reg1<=1'h1;
else scoreboard_00157922_reg1<=scoreboard_00157922_reg1;
end
assign scoreboard_00157922_and=scoreboard_00157922_resOr0&scoreboard_00157922_resOr1&scoreboard_00157922_resOr2;
assign bus_001fcb73_=scoreboard_00157922_and|RESET;
assign scoreboard_00157922_resOr1=or_u462_u0|scoreboard_00157922_reg1;
always @(posedge CLK)
begin
if (bus_001fcb73_)
scoreboard_00157922_reg0<=1'h0;
else if (or_u466_u0)
scoreboard_00157922_reg0<=1'h1;
else scoreboard_00157922_reg0<=scoreboard_00157922_reg0;
end
assign doneCountIm_go_merge=simplePinWrite|simplePinWrite_u250;
assign mux_u510=(and_u1630_u0)?1'h1:1'h0;
assign or_u467_u0=and_u1630_u0|and_u1635_u0;
assign or_u468_u0=and_u1635_u0|and_u1643_u0;
assign mux_u511_u0=(and_u1635_u0)?1'h1:1'h0;
assign or_u469_u0=and_u1616_u0|and_u1643_u0;
assign mux_u512_u0=(and_u1616_u0)?1'h0:1'h1;
assign or_u470_u0=and_u1616_u0|and_u1630_u0;
assign mux_u513_u0=(and_u1616_u0)?1'h1:1'h0;
always @(posedge CLK)
begin
if (and_u1606_u0)
syncEnable_u387<=port_003e9bda_;
end
always @(posedge CLK)
begin
if (and_u1606_u0)
syncEnable_u388_u0<=and_u1607_u0;
end
always @(posedge CLK)
begin
if (and_u1606_u0)
syncEnable_u389_u0<=port_01961eea_;
end
always @(posedge CLK)
begin
if (and_u1606_u0)
syncEnable_u390_u0<=and_u1609_u0;
end
always @(posedge CLK)
begin
if (and_u1606_u0)
syncEnable_u391_u0<=port_0055998f_;
end
always @(posedge CLK)
begin
if (and_u1606_u0)
syncEnable_u392_u0<=port_0012bfe7_;
end
always @(posedge CLK or posedge RESET)
begin
if (RESET)
block_GO_delayed_u46<=1'h0;
else block_GO_delayed_u46<=and_u1606_u0;
end
always @(posedge CLK)
begin
if (and_u1606_u0)
syncEnable_u393_u0<=equals;
end
always @(posedge CLK)
begin
if (reg_0122bb99_u0)
syncEnable_u394_u0<=RESET;
end
assign or_u471_u0=loopControl_u35|reg_0122bb99_u0;
always @(posedge CLK or posedge syncEnable_u394_u0)
begin
if (syncEnable_u394_u0)
loopControl_u35<=1'h0;
else loopControl_u35<=scoreboard_00157922_and;
end
assign or_u472_u0=GO|or_u469_u0;
assign mux_u514_u0=(GO)?1'h1:mux_u512_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_0122bb99_u0<=1'h0;
else reg_0122bb99_u0<=reg_006b4712_u0;
end
assign or_u473_u0=GO|or_u468_u0;
assign mux_u515_u0=(GO)?1'h0:mux_u511_u0;
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_006b4712_u0<=1'h0;
else reg_006b4712_u0<=GO;
end
assign or_u474_u0=GO|or_u467_u0;
assign mux_u516_u0=(GO)?1'h0:mux_u510;
assign or_u475_u0=GO|or_u470_u0;
assign mux_u517_u0=(GO)?1'h0:mux_u513_u0;
assign RESULT=or_u472_u0;
assign RESULT_u1068=mux_u514_u0;
assign RESULT_u1069=or_u475_u0;
assign RESULT_u1070=mux_u517_u0;
assign RESULT_u1071=or_u474_u0;
assign RESULT_u1072=mux_u516_u0;
assign RESULT_u1073=or_u473_u0;
assign RESULT_u1074=mux_u515_u0;
assign RESULT_u1075=simplePinWrite_u251;
assign RESULT_u1076=simplePinWrite_u249;
assign RESULT_u1077=simplePinWrite_u248;
assign RESULT_u1078=doneCountIm_go_merge;
assign RESULT_u1079=simplePinWrite_u247;
assign DONE=1'h0;
endmodule



module output_process_Draw_rectangle_getCenterXY(CLK, RESET, GO, port_002f348e_, port_0163315b_, RESULT, RESULT_u1080, RESULT_u1081, RESULT_u1082, RESULT_u1083, RESULT_u1084, DONE);
input		CLK;
input		RESET;
input		GO;
input	[15:0]	port_002f348e_;
input	[15:0]	port_0163315b_;
output		RESULT;
output	[15:0]	RESULT_u1080;
output		RESULT_u1081;
output	[15:0]	RESULT_u1082;
output		RESULT_u1083;
output		RESULT_u1084;
output		DONE;
wire		simplePinWrite;
wire		simplePinWrite_u252;
reg		reg_00c50bd7_u0=1'h0;
assign simplePinWrite=GO&{1{GO}};
assign simplePinWrite_u252=GO&{1{GO}};
always @(posedge CLK or posedge RESET)
begin
if (RESET)
reg_00c50bd7_u0<=1'h0;
else reg_00c50bd7_u0<=GO;
end
assign RESULT=GO;
assign RESULT_u1080=port_0163315b_;
assign RESULT_u1081=GO;
assign RESULT_u1082=port_002f348e_;
assign RESULT_u1083=simplePinWrite;
assign RESULT_u1084=simplePinWrite_u252;
assign DONE=reg_00c50bd7_u0;
endmodule


